`timescale 1ns / 1ps
 
module tb_binder;

  localparam DIMENSIONS = 10000;
  reg [9999:0] hv1;
  reg [9999:0] hv2;
  wire [9999:0] hvout;
 
  binder #(
    .DIMENSIONS(DIMENSIONS)
  ) 
  u_binder(
      .hv1  (hv1),
      .hv2 (hv2),
      .hvout  (hvout)
  );
 
  initial begin
    $vcdplusfile("tb_binder.vpd");
    $vcdpluson;
    hv1 = 10000'h70e6067d690cfcea9a658e76fdec73a3d4a4cf30ef86c2e471664dc5bae005ee2094dc7e86702b7a4343683fff25271c5dc6c4a12ceed699537e164b68508dab5b2db33ac33829297200bb2a74e49918b5bf89d1e4d69daed193e08772c0dc9655a53e81ee50269cf5820c351e1b6cb660366fab4429e6ca4eb281be4d680fff89771bf1a8f742a9eb946b6557010756af2352ae903357cb09ef4500514d5156e8b0be80b75daabc5e484bba0d382c6da7cade4554cf5ec622194188f38cf718c98f585c06dd92f209fc50702111d5a53fa036bc3af19c35845a8b819af24a8ff70a6ad9be9b5063da8e44a6e8ba0502cdba2667a8f2c2224e1f62fe0adc3a39e2377dbe8b5d66243b7cf7b655a4951fc98938dc3f3eca2dffed9472741ec697a272738aa957c05ca95be2ff9b028dee7ad81d7b9973b0dfbcb87827c65d56c8ab2144c27ab43dc176f69647998d0cce1707f297676b920bdce930790765d1f21b7b9f976cd3de2c996c09f2f3c68dac26097c95a90292e279f78b1a6b4386f80c1136aaacca5fb144c9d697d7cfa38fdec75eebbf6082c23b9dd53a1157bdf762be6f774dffb0e36e8176cdc8a21820fa05043d8fed6a0896c13bc7d3fd0b8abe0a8aec07ff86c98531ed716b41a868a32cb525ec33f4fe2b2212a75189f984d4b23c6d38434f854ed219b069a057338f922f71409dd1c6a0bd818722ed6c426d8c5c9b42757f450d55f082cc376b95b6090f916e571f15845779c06a616d3caa85b3d40397db55c70222a729f7a8cf02bcce8eedcbb118c68225b8be93f50a02b7d43a9af189613097ef915a8b8a3f08a9b189e11ed3ae90b17bfb37c44338f07a720fbba53413839096171ed832a37e4588c559b8d5abdd826e9b3bb44919c37e68ed19203438b706123f51fbb88ca237141f65b5b720b5d0d52743c55adc046e60ab529cff192ece85f7d560cf24787f5a37c655d9d8f3a6d744041ff87f771d92e5fec65313d021c130a34e91413bc27bba788e927762519a9371124bd11f034b9704c01d4664aebe90757e47de3ee74f77e5aed2cc88472895cb8d5856c55fefc49880b5899ddd0cceba3e93cff6302ab57b463637d51afa0a321e412ef4a4e48e0b01b668765d8e8ec5bdb536d7db492c0166c2a89bc00b30121d4b98a9af59048d38b7be37c02e925990b22a52c699b92dc179d62274500df68fdae156bf0e0e44adf3e407d70b69cf1fef3dcd402ba79a622cef1928d4b64d020615ad1b4e68c2c7ba9e343ee061e8ff3ba0e53f1aa33d263a71d3b57ed6f663b789fc07aae261ce39b3691fcec1327a1d1daab267e863a56eef4e37453e04280c943558b6782ba8a2e1170930776f503e4e4d9d6dd792b8c3e0909284e48754bb030b68136536c108b48d26ace766bb38bc74b1084b8a4179fe299001d12f6d15cb780afa52b86b5c81a1c793a4c8fd5f91c947fca27c38246e4912a17cefef4f6d4a8b21ea96abbc971c9e2c2f12b9b8f8eb09258cdd4ca7195dbb64a7876d8febd0e1ad87c163f20834907b69bb3cf7f1bbce77af5f352a1da5571dd621bd1f9f976aaec911faec2088bd277da1ef6c0bc3e903b8c8eda0315ab3859a737e8ddb60592cfa83a82f80f4f14ce2ef6feae8212028fadfacb834a062749aa81053bfef1a334067cbf4705e35593cdcd6d0615269e36f132949b5b25a2207d6e59841a57b766a8f17ac00230b1ca701d01550a7f5974d3f2c8cd43bfd4b7be51f954b095c;
    hv2 = 10000'h3e8948dc0784e834f371248437af0bdfbe2211870f0387fdefac915e22877eee2c3732dbe048cf32ffab0dcdb495d3c3387ef141a0492c86e5a70e925b221ec9dcf661411a919d4a418d7814d60f395767aefd39b2c529b2dec196ae34a27d480684f6cf0258064e76cd6654b237a1624b05f2a29f5fea06d785e52e4d571604df2748e596a89d9d5673865fed497276bfccfcd132c77ec58013cb959da8b159db0bbbced51640aa4d1174be7b3a9f1e878c10f199887fb733f36eb545ddf3fceb5699c19229235002cb144dd09f36da02b0e74cfbee647c95722df744c51df0ead0f6db98344b008767c72a2eff77a057e277f0b320f59a0713ff704f2b2172bc5ce1d85676b8b71172478bdaa5adee56a5b28dbe34def8c6b5c70fe2e91953e86fab3776438bfc4e3f6fbf502927716ba33cdb3f19b6de11161179981b954f17be304c72925801635e76adc46dc3fadc61dbb04b7ce0950b67f837217503e00fbd217afd75416cbc83681a0053d4fe1c6061a493b8f34e7c0cde4b7220b560e9610613bd083947ae6228dc545838e4bb538be6f9d68347aa7bf735747e6ab8dd155fd8b3b3443f3ca970418124927beda81fdca9342c572c2043d795e4544ccc36a24f2594d5dcab8c864c7473b9fc2d3c43c12699760622b5e5e2665f49cce28effdddaa27c3266a561241212544e9a98c1cea35468aa9e9c48a1a09763f905e40a8f999a574c7b7b287ef692d0758f2feb4ff46320e26d55a1fd58c3a80f8dfa71f0359742e707f7242dfed497809492cd8962faafba3174cc47086774885db86d6516f1ad1b8a8f5dbff3851bdb10b672aa2073fd9ca5b5bdcc829871463d8190f8b61264c0b00f8bcae306ba3adfe9e85759e88cf53ecd0e25faab9e827f7ea70fe70bea91531d960983d6bafcc5434899ed1240f26dc18c3cfd19ed73152d395bdb2a09557864ce90de174a635ec428aa9b371d11a209a55d7f74a22afa71b621206a033bdc460ad5d0baf1a6b677ae2648d503624ae24912d53aae0ef1b8a5e12c4eebb96694b7ed2804f7fd052c8cc0de1367b11ceb0784f225cdef16b1eb00fb6a4efc51a39324fd4a274cfda1a235930017f42c8a375c01d81f4b8a92d546f5c282760d8ffcdd9fadc9e97e99db2d0d1ce448afd59aaf6efe4da1ec1482f327232dc57c2fef788a01286d8c0684f176b93a0aba7a531bf07e6a850bcfe1faa8475fbba4b4610b7060949fc452c4dc17f2782687516248cb4593e7eed881728775694317b9e883515b27666283785a40edc520ad966b415fdb76a46778d6750a76fff124345942737a1c2cbb16bbcb4a9d4c925988f0cf91e348eb6e49c7db5d1da7db1f1f8ac9ab71fd043df3199d8d48193eff1d4a450dabb5d1685e3d3aaa99d2a0ae6bacdf985bbe88f7043c13878ed220450cfd377707401ff77603faf7125f36d0951171fd2930ae70aa8bd79401e8b187d0465340cdeac1b94226ad6b348b3b2ca6b18392dc16de89aecb050fa03e2c7615e066cfef89125c7d3eb01e6396143a09edb66c730fa9156961e4e23368d6ada482a1c31516f4663017f6cb9ad0fe2a0dd46e367d3ac14b3d6cb1a39a1495379f877552be4f7e20011eb8cfb8cf7acb926251c4c96ab8c36cc883ff32dde33d4600c282c25527787c15f0edf7e2b446c460ee5f882826d5016b1f2901598d29e4be7b6c4a40709131c87469e10c031e621ccbaa91ae262244a67932d48f4d384ad4a9ded51d831fb1;
    #200
    $finish;
  end
endmodule