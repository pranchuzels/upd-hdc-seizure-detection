`timescale 1ns / 1ps
module item_mem_2 ( // Line length
    c,
    spv,
    spi,
    ch_hv,
    spv_hv,
    spi_hv
    
);
    // General params
    localparam DIMENSIONS = 10000;

    // Channel params
    localparam NUM_CHS = 17;
    localparam CH_0 = 10000'h385ece781dc2bccbd165b943df9f6c66b342c66c2874ae514e0711f121c41f048801feea276873b287bd12f502941a94be1d5f096e25de5e8302869cf77bcd54cfd2d567c57009926b1e29ed122d3749a60ab4bacd37df3243211580480e608ec4e592429b0d1813ab99ea6aaf8c41c9d8ea9896e3baa370797ae8d60df7548c8efd8b349e70a8f730fdd5dbcd3ad80b195b0f7f19e49b9b6f3e20e47646a8e58fe927df1657183795426abe022894cdb1daea13b3b99845b8afb3e1f1407726da678ac5c0ad293ae4e05310e3ac2644596229882bf2a82c245403f0455dc8f76221abc85017edbf8e6d80436a5e61720a508e898697c6c2371d93b814a47c951e2dec4303c93423ce01c98ee41dd2a4fb1c7aaab4b4d7299dadd878b12f5bfc13c678ee0e0fec598724458c4cee8ab604e6828dc8e6d1f85372eed8d4ba402d196f4368944920e7a63def7e41dcfe0092677015d46d86c0264773da4a6d95164463f269523de81cd138fa44eb0c8b34d85eb9c2ecb62b980df64db4c6d6c499e47e932120b560720c0c303a795f358d219c2f362f5842c82a4d0e7dd6616df658586a7bd36fcd4588f7a6e4c727ab29a4c0f556419cb09cf017d1b38a5ea1239deace676ca5006c560972b06e57e58de941c825c297bf2a3bd331359a5390ceff91eecad9b4ed94268b4e7c8720b0bdabddf6a2df752b5e7779e38e12237c5405a945924b4bce6c4a9467c404711fc0c19373d8197ba1906841c9b0896dc6a178eaa81d4d5133b81ddbc2ac9d40230a1a8811990fbcab100b6b72f4d6c94d08d19d448959c65fc6475b59d05cf26e5acd5a557cc0efedea97911be44212482a6d6e1a2987088b49f41e3fcf5c209fc853a5fa2153aaabd682e385e150cd2a78727f8f24f5f2ab1d9bcb2594f4e95c7cf8603bd6f949aed4681af2ad2b6dbbdaa89f1679fe2c537d6594aadc79e8cc290a26bfed7f04ec4ddb84bd40c2372505498ac3d934173f743609de47986694d55948631d0d1bbdd8f6b288d7ca700acd43acf58fc624b570d466cdeae3a122aed1bc37ccd1d567752c1816209087fa33e50fbb9ce25bfa46d9e34eb1386a9637eb0af876693df8540f115b9ebaa9dc012e02733d22d95d998063bafe9dd3a635119757aabbe3cf50961cd7b19d52c59371c42f05b08f45286269f16160c40236958d5868a30e6535bd87311e1afc8539aa8cae1d95b9888ae9f2cdebcb6cfc0feddff96a5219bbc47c5e5dca1e9af4e8119c3c0c4195a842dd5f6bcdca5e37b62632793825647268aafd8ec1fa701a7ed21cf8afba98b9cd098a736224f847f5e93cb4ad107f0f7703fd0b874c85ab21521c252b547e8536c088fee4d0f546c27b1b11cf9a2017ceb49d2b9e0ac7e77c7d57ff196b583de38de2800062a756b9efa9f77a965372c1e839d9d3324d58b4d99c5b89fa9b4ed07103b64b9d49e80f9c9f1da2349c687640f0b87ef32fcd8c6edf32c7c543111b3050fe354b56208519a716dc50d9067a6d6029bfd0f4caaad96a556054fcbd3c5cafff94b994857a12b01ca005581a8627db4cd1df99e1956b49fba3ed806438f7793bb3d54373b00510ca2c2cae760c6dfa93e30725e875cab55af1d49ba3ee5e04fcba7ff9557c50ede5002327bf8e82a1a4d1437f0db183c03a2b52360fbb0a836846cde80f3bbaa656ae915e4cd3fbf4b2bda347ad5b0adbffd13404e1075118e9b6de13563aa895fbcef2f3318c416d0441b671565321be;
    localparam CH_1 = 10000'h45a652e6f1f62085c38a1068a0973c1d214c8ebb67b121a29ca7c6500ff5ec5a851b9f88e88bc2289d420cac4e16871b01d3aad00d86fd14e51f7e26e1239bb261ceb7e16a2b057e758498245d1062b756ff137fe58342911544edfee2674f09f4f1b335c6119ed37b3bcf3af326a513c834609a104e9df40655bd6dc39706c8cdfbc35231292e198b0711045f03a4752f14368c67bf594b49f4d24c90746efccb7b751221b2275ae8c6afda489a147edc06b3b593d5cf09aff8b3e9d90145e70bfadea19f7e8993854d2f542c0f1f25dd5ce4320db494dae5d4851246fa497992fe4105429e997c07357bf6e2a914c207d113fbd84b335b65549a0459a94e2faa941506e6602ba0ec906811476f1aff404d124c79a8e42945af7a65f6ff9fd3001f52089603ed6dc4e440a1df824e0dd63cb90e1427f92b3ecdb65b9bcddc8eb93d2b5a753c06a50ed2fd1617089981af4c6da9a76c22e232bd14a0ba2509f49b68adce7d49fa8ca3aedec474b057b012b9cbf0ea6760f1e7138ed3854504092fd4b483ee3ac98a4c251044d9565f3066f68d81b073883935d3e01d73dfc5f331d585a6ba452f86a01cd9b3cf00cde72408711d001efb953885b02c9dfb0657a10b2b80d9c67cd784212e05ff27467d8f13bc843325cf3f34a59b78d1b99d2d9e132839e5e7ae42840444a5e58a994a617e7bd87d4490db618e865285daa752741aecf45db2ef3a7f953c8afba64e9d97147fc3fc2fd2a010ced24480d3c0318dac14574722aea4696ffb54ea05dbd89f63a8b41440fe30462b0b6a3ce99d2a528f5f046982650e67c0ef929121567467f22b53415ffe4633a87cdfcea914a428db24aa86957d04fec6ae1abd61dced3d402dad536a58630a983ee2c961c7cddc6e1c0d568f804546cf82294a150768b2b013095421ca59cf40b2f650c5bb85cd90c5f6a7097a06d0163fae5a7abb3cd497321fc0742e33b78f848e29fe3b208f932a605d819dcc5d3c09196453512c8228fde8ec85d3d568e5d597e93e572066567d4b717a8e679822027c7f592fcf8c722b6c7e6db2b4bfc9a4e22cee49db6bcf6a72fe8e292f037bafe5e481998b1dfc916b7969b781baef5552c8c6aceaced2c7a188a8136972e7febd451dc85a0edb0d04fc9a2239e05d0813c62066eca3f0ef4ffb36bf17d30ec1ef4eafb60a1cf9f7decd2bbebd8ef00c70950c547e555f02dff66e32a79f372688d4c8b04d9b84e7f4fc3d580482d60a753970e47303dc1e46457548b570fc792834c9d583727e509795eb656f68b37486a2c6b53d74ed183e0506ee7999c2f29771dc6fc5e0da7a72051ec5237e264985225a1da1be5fa0455c257ba308e2b124e6910c1cc2382b4044ec38dda78b74b6829d21be362ea81f2f8fd58f63a1f409d37d99d56306a9fbdcac571eb1cb4b5927f8df121fdc7886ac3adeb43db5f2df50bd4ed41287ff682e0fa93405672983ca4b579d3cfad7a8bdbec5af5857f11a3351ab82aa621a31b9e44b61526fbd27250639c88a1ff0fa86c8092ff2f243beb1bff107d5e4324e27fd5c2be680fbd79094ac4df249242a9beab3df45f4db83117c8ef5c296cce5647f64b17ea4dea3cd21dfd906f18168acf85a93e8fa41ba8b0e790989147e688a0199b0bd4352165295f585560c59698843dba92e48d870a4645c0d9bfb00a5983ceba81a2d5dd3459063a9b5694feccac6671b6cdcd6954fb32069352b7896f589aa8931eb4ed00d8382cb33fa;
    localparam CH_2 = 10000'h442f2f822be27d4b0152c0cbd3c0f8fedea00e23b2088e8cc499ccfa96d8dd99de54d5a58e3c020756ffb05e1d99cc11f75ddff12bff3d9cb6b61d06aa72b904a7d65f8e92ae1c89cc5cb46f502ef2ccf343a548ff5f7cb6b950b2294871aad0e3e36e9cceeadbe23ff97c6c7e0a43939f0d8913191cb28ccc0858bd424ee622908a6b1414071bfe434b82dd73b221d410702f2657a8ffb581fbdc55ad0b411a59aa537fcda1786bfbecbf5da02c1e37a8966c021bb1f78e823ba91736572ef79411c439769cebfbf813d580d52f09a0afd3dbc01ea2b97d2bbf79105339e00d4c7f9890c2aeb7e90bcbbd31dfcee153a49a64b7a3e88a046a2ef774e3de5c8cb6bd8cea307fe142155f8140b779f48ba11b11fe0301add504a93b97ca731d12899a359191d8b44c0a966fd6a57551a151f5cdd34e4c0322984865da72d984743f6c6429016fdbab3ce45101525c043e82727840416ea915b916a4dea9f7709630ac4ed23cefab697b7a5731aaa766be484bd6c32e94e25866a969c52a14588ff3912b55c62ee5d9e0e23b63ee14f05d515142aaddb04e3e27402389d8eddbb0c6ec5d6e477e184d9955268fef233e38b0f474dcee595fd8d281dad0eb96f6317d0b0fb62cdd3708667d1a4b42da8b6263e12196502f7adba6d46c665b6351644c4eff54bea76c68d13492c858d633423ead22886b525e6e75805ad7ec3222e49f76cf953a18205b16535dba26c8d62abdbcb64d295ef982ee080af1a86ab8389298035e9a5528aafadb040b8b72df951447c79226804be05367f65c9942fc532172c4b6b3e9f06dd768171e84c3d2c890a83cc3b935535d48729922e5b931f432f0d94ae2e8af18e5cd172a8a2c2fa4d04bb1645c764e70ca901e814d3ac1be7403f89600b059adce7a5683c4dcac041b7a57ddb52678ad9577383404ece94f7fa195f36cd99f0889e93b00cd75eaced2f08733ad4006adbbeacc7a26c5e66e1f33afd42470f5257c1f289d6656e813ad0f9a8d18f5b6ce6ea44c814c46e20d57695f4a9436eaf2a5afa6a1f72c62df98257f79588213226e978f095f49f02e682726748c98edb4d0661ebf52852d77a2538eb0d2615ea63bc727e1aaa0df0e41dcf0826c977fd116b4a466f676a02372c75abb506c1efb8845857f9a4a6b1dc21c11f45431c07aa69d8fdad0348e0e785c8b5acee8517ce589d3723e785a6b80d00cd15dd880976c15ca1b58a8dff30262bdd84d9b4c0c688b0b4d510565b83235bfa78574a5c50ade58b552fae0ff616b486b53e6c2d44b34e3b2ce3ea977db870c9f8759dd22cd99950752cf2b8c229be82325b75fc4dec129afcc0960656cfd561f1142ef2e16c76b807505eaf4de4fadc0d268efa642e0f86f3dafc939617d103e2d99419703b48d4a74b96a5886e40474beca5874664f2492865c39550ff8c1133c81636cd9cecef5c92490e1b12756c0581bcf4e1a71be4dd30d64b743d2645d842d6c6b8b6448eb51162c776c47d59f471a20a3fa69a7361458f20087ebdc94de676e717687642fe7f59933164cec0aa787d33e5fda595e2e325ab733bd04dda238a6bc050e31372064054be58f1a323a1179839be0eb1cbbfe750cd5916f3c9e8ec80109dc9ece57aeecee21660404a8e3e334fd212d950ad548442b0b412888df9820b552066c2aacfb8af2db50ac2a5e4159d1b7c92e318b33de233179fe682e8511ad6a30550b5c3caae9eef5566519d302b7fe578fc77fd74794e5;
    localparam CH_3 = 10000'h93a5e7159b48e7c00b8c058f5d0a5126698db08eac4bcdf54592ca294cf8f9d2971deec7cbba924975526e735151bbc38ec00aff6c8dedebb80d7fe28aba5aea606c591474738624156b5e73389873d2a6c7165d5b9b1a4c0f01053d91217a419be5e8d44f2125a126be65d3452bc37f0b486dee87e3c11503951f403cf4b20324248fe215f85abcec27307c9a4c1b71a8a8c5242d3612a1e85fec57e9e003601e74e924166e75e66b87b930377f348480e1a9499e37aa9af603aa325e59a5f8ede54d1273f221a0185eb96dff176094370ebdf42c21caef57ba687d45003fc0e253283a956bbc3cb059b149d4f8cd670e6992ceef3575330e6aa798910dc4e21c38ef0800f5eab4f8c2d337f0022dea6e26df4ae386b4eb0f17cfedaae990e4524a8eb7dfe42affa48eae566118977a7d7ce42cc68ba126d49b97cee4ffcc6d0a5927fec68a534b1294e02b97e2f68f9eee3c365aac4b648b3711f8e272612df1b286ccde60321c070cf0ff2aa493ed6b916690dc16ba5392eb666d32bf653e1aab26809c992a082439ae69e0f1fb4dd9eb4e05d3f475fa6641ffa65a3843cdece485a386dfba9982c38f562f21d73e1df00e9b0ad5099bed7dbe1c185139dc1f23e9fb7a2f51f22d1ab68081d92415a460df36b87647cc85cfd37bd5972155025a68d82a032b66cddb8315b3f7526303c5897a45be1f2cfeb096d50b72333f52c21f6a6826275f365fb09e9bd6f2ed567a97b6e243b68381c9446c337587f436544d93c4d83e7c5f2b4d9460ad799372d3cb957a80f436e53fc179e9ca6ed1280b34cfde484bcc62bd13e4319d4248cba61107920ffe12383391c899747c2f4e176b409d409739720e842229b5068b0a797261b9a3fd3df27cef36c3c600675db69bbf9ec6f2730b1951d88f20501deccb873ca0d7c4873d3e5f991cb3154fe0b2834ee0b1a4773f64e9205706fe554997aefd9a9d7d475adf9674970f60d7b4f4810e04f5e64e529e8736f3b6527298048510274dd9eee740ba3859ebf6de0e616bff6664efbc060b61959d76248f7dd8f5c5f7db713fe17efaa094afc24bc2aa65e9aa148c1a5207701ab2df7fecfac337548b9b1eea930e31d76bd9bd3d31fc82ba9bcc5faedcf19b72eddb61af20a7367205f5e034d538f1d1b94c89fdca5498a526252d1599f0dc66d286424c086a1403cb225ea46ca608630c6cf5a1841f5efaf2e024b84847a00d24bd3e58535aef49354c0dd011841fa035dc973fcb5f6d600acfc5055b5b5c9bdb7e60dfa2fb887689c90cc22954ab8582429d51772a44ee68a1f254782fe65c12973b0b956da92cf716ca17ff71d5306b9b27f5664354ef52059ae4544e651273a349914875f0fc4600d1548efb069e8dbbee8a5e95a564ee81aef6b2da9de64712c4a40306fd169129d70b4ef51403b2620a15fd917d79ba92a686b4744d8d45ede078876a975bc395a4382b25c3f5445ab8b30c23422382f29f951d0729f1917607b8b4ba1d82c628712c8876baf0c48c811bd42a700e85524712dc47badbfef6812acd734ea5de72f4b7106e22c23076579ad03ea13061a4cb7ffbc9bfb0c97d8c9894f82e6dd5ea32d642d653300eb85d9e010b228d2f216cb5131e6abde6fa52beb2a9fbc0157b24d57cca7353d954c39aa3a7b69132509675f9df51a272acf4574d58f022084c2a4907143223c4129b55a2a28f7f8250822e2409127690483ec265c18332e0653bd99a58827cbc8b8544cb8;
    localparam CH_4 = 10000'hbcde0061e457d522a8f2e2ed66c59875629f249992ba17e1f23de55dc0c9dbee1d56f650506adf762cd09957f1a19607732987312c648390b38337be41f6c6cd79df8d20efcc044db7c625118e3a3c835517288b1053b6fa1d777b4d2b0e06ddd5d96f36c7bc63bb89b30ccad0ed89531ca9e649612a2189473b29dad43955ba8159ba016163b10e7a7e911f120553556fc534816686d61c01408a3492979c99b5d4adba2ce8fbbacc1dcb17cc948f405dfa8d1e23c6585cb0376be5fdaa13d18183037c14b157bbbc29908d9e976e1cc4ef62ba50431537b7a593c0a5d890ca240290ae1809694b8797904bc334944aa4de90423e6416e9a592bffd476781e7a8d21f96c539cee1c275ff0fb054097a1c07882535fe7c19b799cd51f96c346fad1305c19e6894f89ebe081f898dc7f7adc0942a48d9856478686c04f70ff6f8cdbfda09fa5b6225a5ca7c2aab42579647064ea8cb097d1dd7c40136b61a85dce130bb402f83eceb7e90b15210446a8fa0dd620f7dd59bb868f1c37ec5026f89087acac8ff07f74b1d4d043cd45e9ff3f5776cc10e88e8eb4f2d34bc7a50ef6c4caf571a8a96c656447b72a511f950b6e84f4506088e32105cbf98b59bd6b0bda0dda2eb5bda5d0972482589233dc1d5b13ccf235c7b3b48601382487badef8a3cd81a377d58d49f35481bf9544a04a284c61a5a110610b5b8a185494f547661c4536d244bcf2d528f0a1a71538cb218e047e0cbbe5a6f7ef31b2ebbc5af906e087a039f460b3a9bdd5ddfce96991e0f31121be83771107f7995009a9b63eac04840cdf48bc060c756dd8b41be94c40a1b8fc935765c5aac479a9f9b08c9440260da98b088ba031f59bbf138df32480366b1ff6a76e1690d180e268fcde0305774082f18319c50cdbfa0c25a17522c258b99bdfc0aa788515b30def9b1835ff9bd34017b406c42ee28cca9c2b2e5063b65043dd8ef38901fc201b948535837e872e047b19ec75ed8baca32448cea3be576b072f03befff3c8fc98f1e7f04cc174bab2187fb8bfd284115277253bdaa262f1b523f4610d963de62c68c86c9d57ba78b60b8abf6793f4cde7fbd2912da53918c573ff643ff187883062c322f1cd8b4b575fb0d3df6f61a0743579ffd8ef46f60b5525c28d032802a19c9c7b56131c1050931c3f2a9942eea1180fbd0e2f6897da478fa0964815254ce589cef841081b56288c33a09ed6d2e42145a4ef7be3281ac952a206687ced4a2bbba52bc7150ff5196ccf5530363cf2c5b86c62a930b391cf8ccfd9344038157cd106d2524397515755ac5940f8128933f05caae043fde4597904a4ae9eedc61e794c827adf8afef861fd7b16e90869992c984eac1fcdfd56ba7e243b8a7aedc0cbef981d782089778878e91cd563939b0f8a3e4afbb2038b17cde4b54ca70aec942511aa0355ec1bb1a73f94433bf943746b1614cdb591aead61f46a40c3f4667fbbe770b1cde0cf457f91bb98ed47f002f2d4929ac0a89dbe08de3d4be704a1d679e0d98b005f252cedae6b3a546d0006268c4ca1ed8591cd8a898ae13fd153cf7be696e9bf74c39336fb3082adf5ee0816ec7d858c647139270b0feef1ebedd3b4fce88e476f44ef29d98f05917afb5c801f8f75ac50bd200f0c7cbf5a34d860f197966a2a1c6d7ff29b8757672ea2a23e5bf7b52faf2713a098db27a8d7dc5bbe63b38373a286837d3b7ff66fc5001dcfe7bf647b7b6821578c8e8f47cba973bf49742d017;
    localparam CH_5 = 10000'hf50038760b60d1202db22781e2ff66f297c84d77fbe6c9c8a697e7ed468018a21efd1b18fa52cd6fe13208ce8796414a0b9fec3568c86a7ee43e37f7de778cd7f9bdb63a4a70300661afd26a2ce4aba8259cf7565f50172cc52d7c0e677468f790900ef439d00359696258d504ef7ab89361f2bdb02060dac6c96c672db15c2e970cc7e581643cbfbec5c4f9cb6d3ddd165d8c4592243a1f16af07b1bc9c202dac713337828dd3afec76425385a2426e33fe5df5efd66e06faaa615007c0ef3737c087253e979b6c33450b3af8d697624b396a4d9a41dfc65ba838b2092c9e31fd43b2a2beb0ac6d0c39b435b417cc2a0ff432eb06d13c3fb5fb9b5df4fd1f26c30c1f68da054e116c5de807fc7fd56c920e6cb9b20397f73ba5318c756d717740183181067a3fba75596fffe9a9371d545b79f84f1e706e785b8479888cb970eec3fc8b6148d725e4613b5bee63d9042a1a81dbd3f4634b77c9d740a2987751e124d87b7aea6d554011d47a0af47758280560e2fe25c3a6ba699eea102cfae8881097ff76e98954eb55738be55f2d20b219529b1da4768b2025a5981947224e18680df52674c076ce7d6f6eeedf4c33e49f4df7961bde8d8fbbf035158c84e4f4cd3c840b956f28cf63d68c602f8ba928fd8429dc5e88f5824fe46e45add383febafb4629f7358fdb9c3d505ccd52c0ab30703e523fcb35330afc787f5659804767fa1147f6efab365b232441bb44e24dc8f1716fd47c1432e03dc87a568fc279e154109c6de152543110f6f7b67faac9e025714a997be9c6a60866363115c9c4ab01b15d626cce415713b6e5514afd5c760be5f02634df96e8cdb8d5768acd909c95a824fa971833c75451b1cc69651ad00ba6ed4f43ed12b8faf4ede1ababe57717cf524d6888b71ce4ce5566df2689bad812b0c0c061f538630bac1a752c7c19c2377c6c833ebc00827f0fd1ddb5e4708a678fe6a3b849d3f1572d20907a3f023da40c55284b095fd8b5e022fcfc14e042f67f133456482cf0d0961d1b2a5d24e6e823b313a16183b5de4eff2877ed4dbf7fc8932f4f9343089ef90269e3b20dbfac8cf54f6a89f97234d4dca2b14cf8ea19c1464e5feb181e0f4edf335c2e93e91a8383b4bc20c18f232009cac541011a2acfe34d3cfdddeda77c219e8c8a33ae50fc501f7544a79c1250d6f21d242278d3191eb026bd211da6a95f55426531741986f784382f35b1b362fdd5878bcc1583fee1a39843dd2e9833251470b1c151a5b8a8c597fd998e622dec1f4f61e8e6d60a5ea7f9ad40ba1596ad4616339f21d6b136b80a2f81ddb3f5b8f925f08dce9ba184c96236c6b7882ad3baaaf5d8d3dd2db2e32484049611f65081fec3769c0490bc5fd80fe7edb48de03ad29260b06601600775132574cc2008a49bbbc0298f914a3ef6dd36891a54ed60091cdfe29718afba7ee3c83efb571af3f1ddf9eb967e2349830be328f1cec4622347e9502177462b79e49b7b524c8b46bb2308ec3fa9c0f3edae476fd6ea8c16b5b620f43a9bf6aaea1c00c44a536f3e51a93c1f1d19d15630625943767429d8489db1ab855fbb12d701ac4b589f8c7dd15d18d004b9e9e48945efe2200c195bcdc8128ee19392b13398492dd9b36afa03c3bc7d210426715c5adb9535a015518608b85dff4078fbb536700a1527bf0c87a41c8f6c6f1e2b016630cc490063e64be2cdd301d17635a2078174bc52304a2494dc009ce76253b44375635234879046d1cf;
    localparam CH_6 = 10000'ha5f586be4a6a29f0e6377700a5b10f090b1f169d0044a5210290ec61f974dd010062864385aa2e77b28c5c20e83c84271d3a8ad2de9fe75905141db639bcd653e154d1e1bd2a79485e74ec1f18fed205528be009a4c1fa810edf640cb8fb51b547543c8f306975347be4e0ff06607d856dc0ed40073701379aaeadd4887db7084746d7c60ff50ef5927a28dc95d308c0a3c7b4cf99803c5cebfa930c63aac9475defceffdaaec305affef378a49d11727e0a2a9609f1bb92e056f297681918f4277af43533da73f484f8cb44a03f19fd1f398ce1e933400ee771e7ca9197c5cd5ca9ea192c3a2ea51fe135402929b8025931c101e170dd3ab84217e67be0bafe97de3df9b38622e2d43dbfda51fe77e81e12a132a8a0278bbe350e633423823e28bacf0b205749aed4d58251ce0bb1641f162a37633ef9f686bd567f81763b68d7c13098458dc0892a2c02bdde02ab1b4e16b97b66102dff3a83e241ad544ca7860e62f54a7eda7a7ba891dc4becd5c6030a7407d944af1864207731ea12a2580d362b6e5080824dc314c1d0f9d7b587cc19d867a5d7b43476ab78eaee6b6048436c51042d728ad63abfe130dbd79ecdea513fa8ffc243b6374e442d796b80b311526e06ac41ff896640d61912aab9cd556557441497129fba6de991f9d76af1b4b307a6cf67ecf8219ea8b9db87d889abe63dbea6509cdcbbcc872bfcfc0c1109ac3797762d37d5c8dd8e86545c3a651bdb2b083e71ff98d19fc80b5f539c86bd0c0c4ac16e59434c14b04b21aeafc7021033deddd7d7486cb8e3940ae59e4ffcd24dce3fcfe40c960d7f4340c0e5fdfc9c3168515161de9891a18abb81a5b19b555d2b50223437fe964d4f4c42861dd0ab1f576513b2278f32f1af5c76cc40bd91800fff266e0f4d877068f4917cdabd27446703b8f7885786eaedfa18d052bb0c92bf675502cdb4935ef453ee8ee1a3a8a2358c665ed898f8b8af0c751e76753fe31dd2ee464b8baf747a1a6e039cfe6d9c1fd14a00bb01a4b34aecd90b7932e7f206cf51aea631043f8b54aa83f6b90aeefc85e026dc3ad92382d12ee290dd992d542cc0408d6af980ed10c9b5555e954fc7fda29236dd54e96a8be23ea1f4816b885b8f4b019d7302e5a3b895b7a11b92af38e5ca50ed301a12b295ee2998aff656ed25084b132704bbaa71ca9cb1172d59b19de4a222c93fd833bf907bc088bf876bfa66b7f129b88e9e442cd3431f7692d1381cb129867584fc36fb4d3e26d8d6f4e6d52078ca04d6cb96ae81e413a86478394cfea177be0fa6031307ca7d89204bddc3dc18402b59fa2ad179f0222f3bc361744911efe91ed5bbeca8c0e4185c1243eb5e5f302b17a7243f726489d3a747319cedb534234fb3161fa13055fb00a4772e9b370a9a0917e5538a5d950f2d01c6e543b41797853448fa1f9dac74f7f6d3a4d9067efa6e9e4612d8a759cc01161de1b5ddf4b0739fabe27a715944fc16592a7c5b6d5eb15ad616505e28c6b4e6b94c89278f8d45446fc47ec40809c0da9ea5fee745cc5b57b6f282c14d5d2953792a43a99929cdca75b53722356db0b49562a9a52cd3806b8b98746ed0afd893e5a95b734e1b195545c614b6db78de8586f0282f09de607c723e32aa980bcc542c5f01e678cf7957bd0cd4c576609795b20e4f4f4095b9bde215523c7be2ae5dce34433e45896a88464a165c584fbca6350cafda1b8b45c58fe75ba446056dd5ef5e49af2a43d2b162db4c3863;
    localparam CH_7 = 10000'h14045fba66beb079cda03d4dd9571afa48eb2904dba52c121f5bee66907aa7d7938393de0d7ad453711e881fb73a65520b1e130db95a99dab4a017f9d9df971d4c492b73d08d80e7e476402ea71942d55b6f35676de3103fe7613d3ec350e740668640e6d8d39bc6c2cbf45319ee859f80559cb1ebe504b7e2c289b4360369a0febc6f148d54a067c56d55546ffdd3a7ef0ea13ee0a47e341e37dc05ae041ddf0a04638de9232f20757ecaf8edbae10c910cdc6e4f424ad35cc8c180bd1a0afe0b21ed0887dbba233b5d75a867fb73fe43f1bda841a20ddd9173648194a53073e425e62e60eb601e946c8aa0e975995d5504d1e706a613fbd744da6169212954b7268d1817a12d0d21e70c3e9bf334cc0c7f954f6d7732d6bd0f480404a515dcc69973bddcb933c9a8e29b6e28205cfca64eaf27ccc1a877c94b333767f69321c39b80071f9d579078f1a90d56d41d4bdcc07a8a690733e1d00600601495a74fb1250e68b6795b3a7cc984c591996ff688a3bd430050f14e1c337aa73d0302c745eac9207f272ff2f3ee943e2721bcedd9e7938d6019aefafb9e9630876bb1fcf14b9a3ecc577e02dd325e81ecf0b618fb41b20ee8cb9ef6eafd3637de0280881e91897adea4f81e9469b9b3552c224aa4c13ef8aeb9de1d6ff12448e6dcb38b124a1c45ff688d1e27530b13eb7af96bafa294d00b97c18cecaa47974cb3716b972193bd57fa2acf83865a88939394437d1fe560a2de60c78c8a59e1e33695d199eed361eaab079b18538432496f42f490f53eb8c12d59e2aee45eea3abf18b11cd333e092a01a93bfdca84c03bbf7301dfc8dd640b1f7999faaf5156f7c4417ad55b331d2c99508d35156f23472ae83ec08eaa57dc52f7acc2f21aac5c6cba2923128ece7798b45aed46277a9883a24f032e3e415477059efd4ab3d9ddb5ddd7047230e7b9e57b14c302018f181d0d7c622c1af92097a2355196dd915ccba10baee5f93fbf240905c26b04fc157f5228d41e4da4081408e77fd194dde673d567e9e494c0e58cacc8a1e339b53003021a1662bb4e174c50adb4daa20e5688512841b7a67f92b835e904e2e74ac41b6a74776ee2ea75029b8ced9c7149ede7dd0e848e2e45e0fb4215418c26b443abb05cad7ec27e1bf41d0a34920179aed529bafb1e888f0d18c885ddb210abba887fa9e3a7b64b6af3f948694de4d076e606069783b670e5198494e8699a02848370d6280c54a80b6e24ac0cb5ad286ed673e030dfdb6b1ecab5e0e1c78ed9566ae4e4c79451f52f372b34afdc76fda7b8c97562a31327ec8a3baaa9f12fb1a6f6502e10246aca71d18b6c05a83a0570cc2d31f08ad99ea989de2b963b05e3cb78efc2179b66152219826cd6a57e54b11bf74890b27de91b4bf746700cd0b80c2c35a77a95fe0d1209b62442841e738e568c9663343d8eded8078a636e59a0bfb5dc2746620137ed19a1ee0710849a2c6ce8bee77fb4eab4eb10203a63f35aea150035ad32a19cb97b3521f3e8671a774fb529ec0aa9cecbafef2d01f57f1f52b8453cce857f2bb29d2520de5922be99a0c62113a827edba0afefae48db924f1ed385e97573fd29568ab2a8ebf3fefdf1a6690840df34a220609536d180af04cec8c1f6d4a87a78fdf85064a441072fe9fa26e49d1cabf47ac2394bb838af75e356bd4860ec4311c085ebd7c7f6e00bdef79d4f7b4b7608ca8865d85f10b8b06dd1d6899aff74501e496de7b545ee2a0392e45500;
    localparam CH_8 = 10000'h8146ebd508faa9c38569c7bbaba43868bef81c38e4133ed6cef4c94cfe2d99ec1bfdd0bae0ece1495d6718eade57160f31e926c4f6065ba1fee48a611d35bd1d96f989a6b297184915cb8d14318e9782770a327e5f27966e99b1742641806d909209df58e66590fcbc391587e4ef72dbc19e1f6f13501cce4baa6c00ab928d8890af59f0c033c0032805796315ea4d52113d19b7b8c095aa968d298254fb58151fe9f7f7e036e776374213442731b525207a7d725346b6c531db1d75e523ea149c16102380d4e71d1675f94188c552baea10a754d4520440a4506f366bce31026601506b23981a19cb9bf14cf3dddf69e1103b3b5c791f2a57d882ae3bd7f09b8dd1002a8b2f743406cc6c2fd7d2d7ec39cf017e0fe89eadc2caf184dc118475d422c35ef3985d2f8aa536f8f97699673f9ff3f806f5c3a463452fa000f7a21aa592a7555f549c4e6d2ddf63e9f21d7bdd98c2da9dfedd0c0bb0f11fa50173b7135bb3e6143a127a03a76b0570ee3b255eb17937c20826e2e54efc13c9b1b8a24b4c5113da15a3edace96d64f2ecd1fe77e8750a92f6817c4d8870ab5d8fb592020e385e69d31c7fc2584e05b7bbd88ce59c1a8d1a4e17ddf247919fedf0d4e0229d5de445b2f30a5ade4cfabba7f10a0c01ef9a9cdd8207e7ef3eec7361a6c07dc25aad9f4db8b3646f1aa9ef23583ec64af42856813ee0e8bc6594f490d5a82d055b6dc3032d4d2136ce8611f52f9bd462ee04a24b79f0fe4ad38993e06842152ee9dd48700358604674bb06a420e42eefd41c5d4d35f9290485a3a84cb9fffb95412f916c57caf845d337c83d7f617dab616deea6aa6d374e1cdf768b34b1eb5ebf01210377d0111ba594fbcdc21e713e362a73228b5617f1257a5ba4113d29b609569e0e157806721a01f812cff4bdb3959e308812b622f9d1db7af2a2b97b564c5bbdf470963cd2ae20538500fe933ee7e3bfd251a6769c04fec717517c69d9f4cde621f97632437bfe9bf4458b3368b72bd3b383769f3c881cf007e6ddc9b48d14e4ec242b12e2c127b658a89dc9889365eaa8dbf8714738a4150c5e7edbcb52b3673f6ef16c0f9c8b35ca8499992101d34c0a943ac50da7b55fe026b26669bff945f9fcf64800d6fc420d0a506726fc62386604c21f13f903184cb450e6a30740fb5150757e37c1eb4553da2d9200bbe370ae78cb6b754adf591d9d0d2ec49490e0468e331fe89f62cfed64e42cfa67a2197a4f07e7bffdf04c010e59823e33c1cd42c96c368559074e7cb36995f2fe920ee317bd7d2fbd84f9f38d41bd1b02f26a8a20c46e61ac51ef22c5bd1628dcf5c7caca55808d655d8326777016cc6c25c0f803658b3a498e32d8ca02e9e9a9ae9144e13b81f09f2c3adde33f5ab2425835f3f95467fabcf51c187962390e4b9484a065df0a4f40ab0ee58d0b17aacb190749a773535cb83ac44ec21f56c4e0d3e3fb80207252a06a954efa3bd0041d23fce8a3d7c969184a39fa8a1aa367d1f0fa28efeea18d8787cc4e02ad77269954ad3d43befa67925d1c25ffb714aa1152bb1e305165a2b89de9fe9b021d2a97b3fb0574f22f26087fb8d9c435b183d3c095b666a10b001a3681a94aac0499c0b41c57e05b1f4b40991c3b62a426e0cd59d41506cf98f5056edcf8ba7c19d522bc1e7beefe1877bc17aaf8394c9a3d4420d03a4ab253bf1f2e55b35fab9a617d04a69fa000b03eba6e20af3dda92e46037a3e03f2fc868a006125aaabb69d7;
    localparam CH_9 = 10000'hfb51967a1c0efa08326bcd60cf2bdecc2848a8b950f8e8af95220175201eaed7f485f0eb21f89250e4bb317f08771d17c9749d79e009cc94456fa2c4c1c29f504daf999f492faca34d0309f2780411361dcbb80f0c32e96bca394dbae7d8e4c22cb3a49b880e0a9dc2af322f8c1bef4e30538e7c6752a4afbe69e7116fcfeebaa0ce1c700453cf028a86ee96dbeb8f82f6fb50b870da9437c62013f1a78ce4c2bf0a85958f0af75194a8d57b04aac894e71d542ba71104963d2235289ad20e0dab07f8af949716f713c4bd97f298ed12a2735ca5503719b3b9b0b6fb6a34498207cdba36d05fcdc69371371ecfc41c1a073a427734373f758f564b85337bd3d80cfcf01961c3a56b61187379068c5bb4035079ce88196c34564c3185d9fb93e21f4c707a738650fa80d3aa3ab1b9924e341276d3cb3335bfd80cd30616df4e5cca7c80dca9b3b1276e96ac19d724ea4c8dc4cb36e5172fc7de60d3b7235982bcc83eee1158961b90cf033da43afc844791ba274f2c8442792b04dc139016c44a1fde23b2d8cdc2f5eea64c276d34591785d00448a4a95bb48dd90e0d35a07344f21eaf42239e07347e77c6e89c37e921ea6caa8776a3bff903c14a90f48244c8e4b00ce017bf04266a858dc805541ada8f6ab5ecd46acae5e63a5179e0e29329ea9276bc8e8d6ceb910f09a021dca40cc571b1916d8f56ad57bb9d6f0b0c220e1e79b0a7f9e0bdd1f2f75ff5ae054a786a7b77ce983a192e2f762e782909358a185c253539f8ff4394843ce7fbf6bb9224e03fbea351a104dd95e1149bb8b51b7121c753b0f688aee4b131aae958011e9d45e33b95ab57e30801b5e82c2cabd6afd1a39e9d0f3a1fcfb9d10bfae1e4918354affba6630a05d9f80f562d2bd1b3fa3a851e416ac8e3ecdc1fdf7e9a099b304e46e6ed1e3d4fe545a17f62c742b2c1531644ac701d73c47ff53adf9a62b4aa4abeb9440f4c1270562c9d37f950d66c69a90084fd38f21d7ffc25c4059c2f52b761c554130eff516aa24e7edf67fa5263bb52dfd9a93d1caede80714b2be5117ecb03124f8a219cef998435af3f18bcdb11d885690a07814f254cc03d7f4176d98a93fdfd99b65eca79ef92e8fb36b8f656fdabe9c514c07170c41ac6da418011c550bd6f0f7ed9f053f1e35b43fa728723eab71b48b3cb5b70c29867e6354ec63a7aaf73a7aae5df7c0902210af54112d990f51ed58ba6ea201c3d469ed67b76f0ecd97c085093ed69a8aebc16733c3315609763c211d2be4339eb807be08db8cc983bcf288e7cfe792cb3cd00d68ac2df08613f746c5d6c3220d1caad786debb8b7a661d83b7dc93c59f62773631dbe583563c1f29928c698052bb8e7e509558d408e5929e2b7dcd2b88c08981a31ccfa6ce6f4e0e1c3d793abc61be5283fca398015ca1b00f58ac3a752cd1e924022954a4b2e5853f03d5fc58f8c2604be2a9ee3a3c18f9343906fbb14215b9ddb0d98b77d934dc7f6a87ae7905165835b637f3397d50dd9487befb8cff42f3f64019299c42e86588e1092f11148358fac39330c2c951fb9bad26f720b7515df58c167a4ebb369d04f13a9302e8133b664f6755d3aebc56f2425f3643c69f01015b20d582d2f4524784697054bfcdc17911e637bc7fe25ca5ac584889178dc870a107a8aea9ad17bf53136ec32463cc73780245086aa42737ae7b825df6dae608a5171e1cf77bfe84e86ea03cdbc82a34cb46aec300811dc830dca0c0df25d75d741;
    localparam CH_10 = 10000'he229b78f9d0f3832023caf523b1406c78698611a0a62cfafb777e14ee5e27c67983d88fbef42346345519826cbf257fa7479f865a85c5a0a98924c9d39bb6befa83a421b32a4fd6204633f7f407d9bc0abe8e0d65cf499ff80bc526bc3d6427b48ca0e6e231dd335f7eb4c544b8920a177a0a24f8ad0e2c4c9fd6ca401e65f53d2acbb347c01939bd2f62c0b85aaefc86a35e5dabc2f7dbb03c2438ad51ff65bfb66dd4071a1479cd0d88a658ac246f03486bef570a8718b6622d840243a0904e8c2504be0525f44ffa17608a0660faa591308f80c3c6e47eff028100c4b071cfc0d9fed1a1470c32fb0d1e8f0bc47b51aa9e933a9b31864efe81d471cc486b4da0c4b1b23667ae81cafa6f66f239829937beac69e1b9d6e1568bb3c7ce11125b2e1ecebfb6cc63b4ae375c8fb7d5c3844581dbe0765be29008545dd614f893591d45ee4d7964ee081744d300fb29961b14038be330750ec4f47ec4ad5ef34868969560e52c64a154fa0518565bdeae0db7aefa252d56017815a3540508ee3f95d2f49751a64595d292c675fe13cba4d709ca229e3736ac8a9041c5baddbab21ddedb035c90f95d0d5852b025ca4d289cf6792dfe90ec7987397bcadb6ea2de6adf8fb7d7b33d6add768879bbbb2cd2ff71b0acb17fdf36915c60475f9812d17aceb4c4534e3f3590990cc07bff0793a691f846ece22b350881220f75b1d7c6c1258c3a4b7370a9f91b61c0782b39f23c89219edfaa2531efbda9d597d9fbd7eace5f4291b2ae8eb191d82e791e355444c0f8e8826298e57569ac6438c6dcb534b5cdd72cd6a07f192568c7e39e0fcfbd3fdf1a98db0051b14d0050ac9b60e4acaa9ba75eca44f6c9a48fd6d77f00d454de1ab62c31b977e238bd90f79f59730a4e62590d38097fb6359741c00baaf8e4465115b4cf3fe3220985f38b93063c3bb5fb1b2a520b7f18f94c3819bdbaacead5ea6bb8b5aff7b786a874d294337f7cf750af40bef4f39ce606db964722ea6edb974892f3ac3d4e8ea0287fd992acaf0a4f40dc2b5d844abf393f6d3c25b44a93f414e2d4158fc46d2da241bbded4eaa049ef976cc9cdbae27067c54f076262fad1ad93158a2a4502f665a87f918ec9c1346f36dde451dc074369dc5ba97630eb875aae0b66abffcb715ecad59712313ae879c124c77d56c863281956a20fe21ac0b0b22a9bd944c6bab85ab2f2ec8ad02a98d29cb2fd5ea9a1bf57e804ede1c1f504c86e0dc82f3fa70babf4b485ff8c492c8aeef3386cd5bb75188c423477bf17c29197af65497e0c76c163dbbff5f32d568e51a3edbcf374dba2062e85bd6c2015b36f07f418c8708e7381a20977b54dd7c5ff052e694e480839f7ff136588a9905e3341121b476a85f66bc52c370a6f9d553ed8dc9bef20d7302f4e804a874dd94d78c456c111f550e78f49e86c618995156f290389d7ba80dea2681f832808132423002db9b5e0fbf8122709565b1e9d263572dbc5287f4030669195c4ab1111ebd4391df6869b1d4ce45a92fb503df4c906d2688310e9899f9bdf200004aa9a1f3224b414808fbe151566782b61a8a9b23a183c9d9168fa01e550d21efa1abb60da25b6a44e7d1183b932663f1747329fe02269c1284840e64bb5a097e75b85d90f5e0c0d21090e647dfe57d7e06bdbe38a9df03a9f54fd51f58932e43f6c262ae6a7e286c3c7120785a6652abb207f9bd14c91218adc905b1f981902014d00c03ac01b107a82cdd6fa1d23a738a;
    localparam CH_11 = 10000'h4c0334fdc20154ed1958041f37ded872853f73f322a9a1f416f3bfbd0e92582fb0388c44506465440d4baf386a91faf5fe7a70d259261173e38eaf1f3509e820ca1ff087312d4ded08550d3c20289093bc9a3c6bba3fba6817474785fee09dcc46e3566f849fbe475af34cf805efd33fcabc1091f3ed69b1885ef935a554cd012d4de3f3795a625835e857fdff6dc1a0f4840cdd6aed369ec490b78ddc0dbd57fa1d6ed7c03391c5d6b9e17ebfc1e5979ff7a235a082e4a67623aaa22cf01f1c34710370ccece0a82cbde6a39c226b15dc9d6d53d9365b830496965ff613919b645385cd76665b7868fac751505468c7bb7d08284284cc9033c63d853e3f5e14a7c141971d93ef8bf5d240ed12b2426a4b5d3783f87fef832fcb04779ee6a5ba9c12dab86e39216552d2922d9144aa4f47271baba1ba1b9058f4e92674a1102761741b60c2d1e389e4d005ab085613cae54c452574f92ae15ae12051b8d9e4fabb1e385655d1670d7b86a14105e481a4daef5fc0f0609cf486e8f5b18cdc6f117add54e937782baae4279fcf14dbe7d22d09aac39113c413d6511ac47a6965faeae86846fdc0c1a49fd8f884335b3e2ee5525b377b05fac0185b9a2d539a7ebe537b0e793a33f0b68b802897f2f5d32e0a11f9f7a5481ceb91cf0aefc412d7726a6d4f25ac144718c31ef6c58a12b3631b7cfc3d8fdfab59b63e14bf6f17529643c7844b00e7e1affd229c8ac9de7bcf78ba1b6c9881a136a56e7ffffefc9f8424e903c5eba010beb790b1a06137a45c645dda88f9b52151b16c422a440bcbe52e7d9b23905d0304cee2a571596dbf2de82d7c0b50603647a3cf025fd21d63c16305b2fa3019f9632902306fdb4c629ab1d2ffd53eba80ee9489d36bc673c7b74babe29921db403d531efcff37c66e7d5d4b3a580fd0fa26bfe3e18c51b4105a1737935a6919e2c3de15131cce31d23eb1556470c994bbf7e5b4f9ccf55b484700fa80dd1c5ecd77556c68e48cfbd20c591d7fdf556ca83008407e6a22b310c4516d9e7b271cf851b621fac0cd2a010c3e3e6034983adfc1ae0aa58e19af55c7129a890b0cdcf948bfcaafd81759ba75ecdf5a6218c27f4dae604f7d20a3c6b7f43f761672b05dc3b38285b21149574c4c03a947ba9f7a7105036cccb2ac231dd9ec0f0c1e122c0c3ca04ec0de9ee8bfb8f2daf090688341d841a42dba1d65dae13de8644e35dae82337926299fb9896029943658d3d9814962c5d720fef55006ea73e9e45d61f84acce5a0f0f49f7147e058a4735dee80eeae61a78e0e349d65dc463e94589c2d2db2bc76145b5472d2781da2e91c6e4c8c87e14344f062b01d16eec0f7b693011cc4d7b4c3457cf334b349abe9f9e7b4afe840f6cae2129cc89f082bfbeb6972a26afd33701b38c7832de74df091e07c5a773ba7a562c811acabfbc6ee4187ac8d32a41a9f4c12f4d1b2647508d2318894435dc65282c23adf1eec7c40290af8a2d6e69083bd8a52dad7862b6b30a0f0f4863f26aaaf1d7ade94d0e8e9f00db026db764949c56f6f5930c58dbda3ba7059a0948eff842fe19b4fa1c4630a7c83a2b22b4d39721827a747c3e6b27045e5f03769109998318678ef097d18fcac0405080fe331bdb594dbb484208f5cf0bdb2f94a563ce0c4b7a7121ca67e4379340e87245fcf7a5492071318bba41f300f59ce0de37542af39548ea7ae9eedd8d1d69e5d8f5346e16168ac3f2219d8c50fb825a2122b3b2a4153910;
    localparam CH_12 = 10000'h6d3baf1e6079e22811710f54471ea765365d6fb72e00c7144868ef112cdf26df50a500fe43793772568fef1e5fe28285e4f350ecbe503a3547b99fef063df9923043896bf2b435aecfe7e7ca2177f5f55a54b576e6cab541c1cb87aaf5ad36a13cdf787eb42ecca1cfe5cbfbe6b7876e14a65b920b37751cdeacd27d84c7ea67c51be8242907ee2492be389ddccb9e109e9c1faa8f4ada7576fa0aca0dc3c882b4fc8416bf51bc3b0a8a9606bdf56c5008c078e2a2a7680d90a2f6cc3cff1fb4f999fb67431953a8139e8c93aab3be339ddb12b8301b0b068c8836fdf14b7dedf290d92d14562f4e59750ec60a86272a0eefd31debe5940ee62023d55cf8a594ba12bb487977c3b63d034e6658bcf4b4bf24a9b65f70ae49a1019aa16627dec6bdbaf9e4c3bb64fca6d9531a893a031f8b8f2d3c081935ddaca13495de5f07c27daa6e83090f32b1b0ce97af931e5f69b48792690df155cf402ed3001b7bffed00ebfeeaef1ff408c1959e9fe5469e1f2e24e86c5e957a90b2338536193f88237786f4d059aa50cc0304612464a66122e2c0190901fee67fafe112a7569280042565748488fc8fb4dd20a91301a400de1133b381d9fff83fadb3144d45ef6864fda78163ddc10a63c380cae10a7b1c4214fd9e4fab430bfd0bf439a1056b433e5528df0f9236e23f352e4ad7b0821a1388fd3c7ce0d767edd5d41814552219d0e010c7f521faf5796b8e904a19713755b360ebf428bde4c975472c6f889c93b3ecf1d365d010259664f22cc022e820e133a70a100dc88ac3a58a3fafd3e2d3ea0e1b2bc748263501678a90ba73b82044135a9a6d324d0c53cc0413bed9e70402776858c9b9cc48ff5a5f05b8aa031ff1ef1ae45ebf4f08dfb4e748b1f99132defe3f3218da8ac41c5dbd5a716f1349ec773c9e8c6f5c4ca24147e8d71033c5ee8ae55f8ede25f133bbb2191ad8948337dff42ce49473e32ed5b4b52e06cc862176dfc04b77c4bf65ef478f7b6e2f6a7ceceb584c91bb32b430b57483aa173a18cb9f9aca9f0439a60200413b03aa6afa0840eab8cf55178d222fc5014dba9d635313e2a52ed062fe6af978773647a724a87571e841553e14c0d452e1acffbda8ce0d881f130e62f773fed97af2bd6cde6fe53bb072a12bd84af9be8bd6e1a8a0b0625042952d614cea3b8c3608fb952d4156029b951c5a5cc47575bfbb73c6da4799699692731b43e62e347c09da49e36845baaf7ebf4a158249ae6632bb2a005d74ea5b9f19e08184d2130c8b0a173b5adda6114ccd08ebbe51b1f8a4a7741898bf848020eafd3e35822d1092f96733e2304d125356021424bcc194c5d2b47006346d653236aa3f9602a8c04e1c2bc4b82dc7818164145771e82c304fe8d11c7bb632af63c1c2dbe59ac1548c85060f16abc02d623d70fcabecad72bb0071b368e34667d31de8be74793dc5bc7adbd50543ee843d3c38ffabc6d24721acddf4488a10fbd4d6527af59bb33dfc49c4690b5a7d0c425072e6eaa8304f50c512eb895d657160e6b9d30fc051f75a48287c44219e137de5d9de79be42493ce7ae7b99c69084d0865f4c3cabe2bbe4b7849e84507d62c13f5066d4b81861d4cb2c348391309f4a571d37d3a5ca0cffc810b71457d7701dfd16b7796a422e10314e01e9d345077e6ecb6946d32a571846b8c1dcea593942068aeb5a7d97ab3c8cbb2f83378a6d99f5ba6beaab88e9a9be914c55f39e8accffa040de074ff9c197112c0f25;
    localparam CH_13 = 10000'hb17edee21c0499e11c37cd22966142430120a93689de26835f3fd18c88b47f6b9c88dbce673351cffcc43b695a0f9f308093abcd622dddd076e95d3fa8cd497c0908327a6a9c919f2a9dbda426eb511a3cd44500a0b96f2c2bbf4a00b6e6913c05a3a2fe9dc7889319be6e1e7cd0a0cc0164f96d7c82e5d527c29b594309e8f74a052636b8cb07a321bd69b075d20857cbe19d11eb955c101f5a100d20c011c37eb5375face2551f1db309d9bb722079712782f489fa90170aa0debc44737a2d4064724eec03779ce287d9978a2652e54d534fbf840356774fc2d451d874bee062d728ff7d4dbfe5acf75a8ee1964e5b9530ad688806146061cb0ea6fe3abe9376250b368b333b7e9f5b9f208c270d4920eaa5f72aca144746cdcfbf76a76fa4a64d431b86a895fd11e7f8cb9b65e35963b3facec6350f03393e2069004046eb14f7184dace6ad80bb3bb965c2dc7e5d43dc821fcd07c8c0afc7ea81b7ba5ad634c505a98e9f74c3f63fcbcd028fafe4d627bafb16d79195f35a31f13cd2f78dcad11c3d02103cd59752f48c170d7f2c7eb9b94951cd48a59617896186714322a12b71d760d38939e0d82544c45c0d75641c29c0cc031500e10af304d8e00ccc3f99101ebf7d2ea4259760a9e39ec32d02eef92e65c8ba27aa63b14f6cf5fec84593b58b9f3cc0686e67b9c660affa5c90af112fd035fa64f4a97786bc17b588f35873fc64d059d023d2b822ce9e8c1361d2c0a6cdcdfe37b9931067479987aaa11014d8698aa6c7026fb12cd3a90a3f8806c7c6b35dc90c1877e5484e8e4bf9b78126bd04b13cd96a0b2ebd62532c5409f6203cc01a9613960ab5c964e6edbbed3f73e7e7642e5242ebb2a085932d1a7407231dabff2ee6ee89f4d714c8f40ff398fb96d9efa4b2869945468b5f9763a6ce0c0e0c062bece3c126d8cd4b5950960e5ab3d5896e081f314d3c22031d0f9933036fbe2c5ebd0752b2376b81212880ea695dfb613379308d659a080548435c5b64f349d08780e0a463d4d9b244a75e7971abeedad81c8a62da0c6b9324c933315f291eb16985b5dcab1656eaa4b38ecf7b8ac36742f76e7dfff10a89ec864a55de23be714cbab80e7b8af9e857f3974123aabee8679c7a26617f8ed2439c4b428e46051adff1d192c4dbae0b28c6ba45bb2de9b66a46dafb240b32c67961561eb76ad25152c6971bc1e2f8aa724cf8ffcd48023185984085791524904a5fc79da9bc5d58c77061fe816994186409eb61c0aecfae0f627cee56cbe280348436332bd9582cfe869351a979ecb28cfe1d3a56003006b4020ea1ef9c67319622559f3b3250d3d3cd5042a9c51798a9f7b2e2d55265aca8cdba15ade6652c7523a50ed9114d72469ce4a33f64b21d6f6b7f221561211ac363488bdd30453fd3760f323bcc173c2a45a1a78ba6319c6ed67497618cff67b942b24e59837ed4ceb9f03a1d174b10a17b629939c2d554bf1fc299f8709b8573559abe6b3a8a5f171646c44ea6fae271b4544628744bdba98e43b8e45b3e74cb6d4b20160b76bc77bdbe30058aa802a287b5433c90d9ecfbbaa04835b4d4f45af6988a724d905c3f907c62d15af153457da1f56b7cab97fc4e28a5b88d289da30ae5d112d5112ff4fcef657d27f01d682fb30effacedabad14590095f0f75c93dcdb3a2c29edb2c3841abaaefbdf7af95534c67e38d261223f21af93777f76586f4a62c7782d282d563355d48b3b10edec9463cfd5efb539088e2a;
    localparam CH_14 = 10000'h83fcfa39cb394b4df6a609090346e9f401888f0cbde590aac63e105eb6343dd0f8d6ab323b8f42135e797d99f3233b4826c65e51adef9e3cd93beaa152c2e298f9ff2e7aadc4112f77c91817026d2843f78453cab4e963e0c325e2140a55c735a0acec3f9f94c870807860e797d8af1dc668e3e5f23e326ea17589f91fcc51b9bfb6bbb5353e38454ab2b736b7a5f625f45bdc2f430cd7129414d1bb8cbd0608eb3129347e9bc4a92ed1c98dd865941457ecf6e4d7e95f213d1ef88924c954df94cc0daed8e2ced08cdb2e3b386438ffd528cedde9cee54a73fa97198870b9b0a5a9018c095a43a3090605b190897b11ed0c5b985bdc8c080bb82ec5779a74a309c89e9f44ecb241a055bbadd928589f62a22eeed14e09ac1348f99d7236e9b7e648e9323218215dbf9fb4d4940d20e427cfff63ede39a673048230c492bf2485ec8262948df40e187c92ee1eece1c9bf38ab8f6e60cc9ca5a1c60d50a0971b2db4e66a911b9fab06afed28a127ab1d5ab9d97d70ed3abf0e3f0e0b28be0b23778093f40221b32179e8dbc4f69d2435950e587afefe91e9d6c68a9d66c04e90f41668354ba0750517e3f2ac55e65904755bca20e9dc1e9e10d68dd6ddd9ab3a318be0181f430f09308f356f5e3de0151acef8fd7155dc71007a4e14709a9bb1084763d135dd1ac923a28b51d2d59b0e9e69a66495bb5241ad1ba3733dfcd20e4924a69df80d17fc465a2aa6d605ac334bd6ed2765de6373fdd6c34a32bd020988fbf21ce3f0b286af96ea0069c12074ac5a9549584c591c7bf483e36ae99805b7a7cb93135a1c7cbc589ca4a8a9891e7b2da413550936e0e6411238e25a0ca67a71e068a10fa85431d44c622c9611c256b3a5d6e795fb0580fb8a674d5b1d5566c20d0e5ea353f533abb09a1d3b6181a0de237c3fbd753df066e15ca292ad8b580407acd531aed681b2f54b13f9a1e7b26cae3c30ebdf5576f2a9a47d9067f0e420ed32f9f3897b7d10f5822b891e2b06380a0d7c8b29e6a4f817c47df11795bf47aad3d21582c42f55de464516b5d913f61ca08d8b311e9ba97849deb9a22cb9358841bf518f662ac7f7167a4e158236a10eaaac3680082f08bd24907be2a493460531dd015be075fbab77f4a3ec510b9b97642c58eaed86ec33d22500b1b227ce99f7aeb3c5c061db9f03e78570c3dcce2759a0a3f1bfd889bf448a93207643794a96612a102c8bcc93b8c44ea5c18134c7105eef89dcd9ed26ab335a73041e2ab4a6746851a02b82e7d1a3821fdff634f4991ec53b6b5faf7d76779f91e091fea398b0342fe4b59fb51771147ecfbecb57e01d2e3adcac7cca4a9956f4a0afa7a4643c56445406d85c6119460ed74cbe9bc9c80ecfef53d48d6a22100025ddfdfd9802a00fc6fcfa74304a670ebf0c377c3af3678a7c0624d1a5a3181dacfe8925c81855e7d684bc8d553cf0037bedc7d00b6dbcec7dec3abe193cda790bb59ded9fd27852dfc447724d427fa7129a2f47c746146b76048aae672b2ce0b02f21810e30d7b4c8dbce9e5ae427d6417e1d97345272c6ca591cf0117dcd5f2b16a2b02e5a02eab22d28b9d45dc4b8af43c0107c6a09e5993f649bdbdfa62157c931364d7f25a5ddf9d879d8759166b2f126355955de951424c6bd49e0efcb76eff04410174d9b5fa15203ad69e39a6c3b658e8e673de0bb8eb6faf96dd2e2c86d0a1c1848143bc8a384d84abe2d42476a76b18f1fe89a67d4f5293a653d548e2aa05;
    localparam CH_15 = 10000'h7f8d695ba751d1582461e6752cd3260c02ef7a6d8de2ea48eb134eb1517f11635c3a1a5adb04166faaa9a2a0b228f234f9452ae8ba2261833cc2164dea2f90d495e93394777ae6c1a8e7f60efed13afb6cdd7189ba415f73d0a014050ac6979e62f68ac55ab7fa81d123702f0d0a4cedc856cc911efa14c808da645bd8d09ea342a5898d285eba16f96ac8c6c42b2c962d46dc1c65e7f989c162e87290d19a4e10aab095a1bbf25abb5f837901ec4d5549021a4078e2795f2fab4657b634f8e30cb72fae4a3b3740bd031a07e3e7a6e57579ef4174bf5f2c75bdc19d15f5d74ec96827e3f15b6fc3409620873364ae462e9cf61c6365b3bc93da84339ebf9799cee6c50766cd3fd1f56e44df866039df12a9c0e6cb9ad48e1e2175996869f12175cb93e18c956edbb181ba2e412b2258348dfa615b9d80eee0c30f4db72a10917f5d3f1d9ed570e9b8bf2390928b5857418822e6ad65be5063933dff3f9b3f8ced6d842020f175aa82667b0f0f94ec94dc7a4a950adf0baf071caa490bc9007b2d8da6513d8cc0fe677368747fda7c79e159c5ff440783324d52d156d56859820d6daa8fdfae84d53d4beb09b9f043c277158b16077b096f97031c1a5d7940c2d735e226312d089def07f8b46d5d5eaf872da1f5a084078022fc2109840433f555dd4603149762d689635d6f4b1d6d24a48a825986be732894c9bbf9e3d04ff36e73097577da9a437d9aaf59f52ef03025ef65757a97d74d296eac89d3112fa50ca3621a4e1b2ccf35f8fc20cfc521d6050f993b341e2848bec1efb75f8190d5fac3a5948c3a3c8ef4223ac9f327339ba94682b5ca6875711a99d012649d49036f817aeb49fbf349c060cbedda64f0e8b45217b329ab3e3c75a918a22922ed65cbdb1b42f864253eea35a2e0fc690f52578f66b56c1bd31ad05b8c483768329a427aa30ee93dad893c0630aa29e3316dd743845c9123c18400ea80309a6d68378ef3e3c0150f84a3f21fa7d662a8757c48dc2bee28babe1324f7515d226b101c847f33c8fb065dda6efb0665d2b45d2beb11895ddd77194a554bb8a03596a15bc9fa40d4ecea7a772818f441f1d7a94362ebd49959404ee9e615bf3d078f93ec5d1585e2674ba9c029deb6ea8e8cbfad25fbe96c4627e9deeb9e4ec648449c47b15429c5d5546219c8b9268c6327eec261fad6160dc2c63f395b6ac813318740839007c7a755fb06b8c22d7e6bb490190f8c14a3cba006799ed0751f029092361e8beac03397204f0e88e91bf3769aadc936c72d33be6e40f0cbbb1ca617912e809fd928b9b60e58373a11f6af3ff25493b05d6d6931755c407750a7c15ca91442bac06b471bca78c48f2b80f1880718c7d8f26c6bb25a15db37c83ed5ecc5ce589e251f1aae207d1c1f23c5df743cc72e5415b17bb71c60dfc1c46beef540f611d39ab112b0db10ceef23b63f94a2a6b51e696c04c49016da5f45b07248bc44dd89b74bd6b2efd876319943c9ecf12ce3219f210272b16de9a63c75ca70ea6d0d1004b738bf1ef527b428336085e26bbc3cf3f63beadd6d988e4009671aeac928e70dbd0489657b1e363677962318ffec9aff135d5ebb703f0506954dbee3ec8f9d29e16de484ff6425e80e42c2c3c0bf74404c1ee035dea3b9c80a9511978e946a0b32542145e1302002d5354e5cccde5ae95f402a267c2837ce7dd99499e5f90b95cbcd3f9de348c5f64c2d74916ee7bfbdb5f2c714db44c2f00e943b313b63db;
    localparam CH_16 = 10000'ha35deb8708c2adad762d97bee5e36abb501b28064accb6d6327fabb21bfb690129e6419e152cc5125503b9d168da70f2dc7373238a16ee1a22e59efa0a17f8083553b11c23b5da371527a6940298455a2d7404335b17c597d01c5d7a270da87840835bcac88e92753c9d4ccba97e50091d4b6ef0e2c7db717ab751578cda5ff355b74f5354bb9ec274064a027b0587ac664e9038e3f61a70279607ffeb5ca411b956420498337a8e1c2ccc5a1bcadc8192bc55cd8d6d7510655295027acd9c4277a6ef4dbc087d9d5892126e35da7747294d19c7089f6927cc48a6423b7696b98d79b75295e094472fe3df31e1254a4dddf5a3b9fb4e6dcf51d5f30687602370051bf526184086a307fbf2ab76ac06d1848cc72fb275f07c68b3ed33635266f9692128c2e0cd99e82a21ea7a151a260cb7ef34396045691df263c00face42bc9a1346362c14337ae4b379640596c9112530595e6c952a0fa444a8a0a3d90b9135b5c4445d3f41c2e60b884f1555b6dc26e33ddff77dbac722ddeb5d8e5c6a54d6a82f02a98af2f9e6c99e624e2e9b6950a28a04adacc0ba096eab5483681347a07c9cf8be483e54a879b54c14672d8a66e46b133985a72a64e72d526ddcbde22123cf35c900870d5e1803a6db0d4dabb5b39f3f866130c9a944109eb5c9a235ffa99fb915e515695293a1a2c7da1a02abe4cd637c8a2cedb43cc8f7bdaff7ab64a2ec467b7a810d1685e2cdebc1eb3067615b454349ccc6ddf042985e1171fdc28bd76568cacb3e4d0dd459be772b4866e966e2b292cf813556fe00aa11faba4f842f36ff5073fef7fd0485af37fff9bd156bfc343703f6e31bf61225280ef32a779d05ff43267f8cf9bb7e9474a29ec218e673886ff10b7cea78e7e536daa817124c6856a56e042f143e3a3c00a67c7e2d7d9745893808ccbd8898387d52133b9177002f2514d9b767d6943c9cc8a6c325f0bbbaa92a21170ea1c9f53e9214f9708a6cb6a4e3229561a9a11f2ccd4557bcd447b1957535efab3624c3841f5e42086cc55a1c38dd93e14a039ca0349c82b6a1c1d301202dbf38db9b8a3b67e824e2374696235bac232f6d680c6946df6aab3458e659de9235f7f5b908641e1d2e0d693d373fbf3425f66dccbf362433ceaa2c5756b826f5bff6d5b6a336e968305b6ab747d85eb28835624f2bf7c97db64ef986b2a345d6fc6d84f65726ebfcf05a832aab349f145771ecb8568ea05af9919d252a971359c277b9866d262ab05989c398ec19003ee5f5dbfba9b101e85202a457af6c2fe88f1b99a92c692639c532b93e2c38a0fd90d6e7141ca87e434247e8c6abd8f5049daec472d4d91e3538aa75f35e8914320cec78f7a2c12fea56493dec37f84be81a234f41d7c1a022f27f8762af048b8c910ebf2cea93d6abcfc354c44451066fadbab0d97479b840f3524fb612457b4b79d25c11ab93aa1e449db7e7a2599f03ce4cb3e945d3a0006fcaaa304589092183313318761ddc2d1c6451a04505c0fcad640182c9f1758c88c9381150ac453f08c33b16aff26bbbe72403a67a1565a076f57efef51259eff1e72f54cc650d5362ca986d019fe53dfcf4283513e15e48411e992b9b8a99ba79202c447f77f90cf2a979f3a17bb8977e834e29b87e33e615b7f26905a416038bc8ad74c7fa250cb64b9d42688871740119972936073d158e2b77ff65fc5f62bbefd8d9f6e36bf90503a7bdf63d81604aed00d60b8caad9508429ab18cdd1fcf02e3;

    // SP params
    localparam NUM_SPI = 6;
    localparam SPI_0 = 10000'hc7b1f73eef362348e22060bab1862f84ad75b8653cd5d7f1029378ad8814ac2fdabc352fcb490bf3ea6ab2e799830b1c55f000a30ec1b9707ef6b16154fa4514899f7e85a2d4f39ca54e0efd4d1d263aad9281ba1eb965ddc23621001032fd803abc88ef6e7ce12bbda62ec9927776d6b6d7dd9588b51a90b0b9e9e9d8ff06d9e9c0c8404adc8e4f635f98d2b22074f4d564c0a8c0d49d8e222401b46f3f5739cca356eaf2199b67a2345bcf9bbe74e0ba4fed7af8029ecd2a2901150d8216804bcf43a1f5f191804cbf20b33c1c5c3f0f70c63408afd2fb6fce26ff506cd00a795012ecaa2616936962dafe2f2c3256afefa2867b4318480b424983e7817107acc9fb82251837e0afea87c36ad50e7058ffb04c5e703838414ccbbe2342d4c28fae904b6c516d11b72e3147b334683ea3679d97affe8a8365312fdf5f4746ff4080dd50253990aa304a80bfdcf3d6ed985e468c72fcff2d7da9010cc34ce72edf0304c3aa58af0ace8378aace09133107b872662572cc5dcf9e62f7bee3995bd329c1fe60e5105828f222c217c9554fdbcd32a05d84c38ea6a53b1aed87ebf4736a1198a0c41086b29d35e84b5d53af7156be50c31cb3bc65ef839ca72c26c34a6428f3d87f24fc5fb16e952362e9009739a7a2f7dbcb661b96eadfa6bda780fad271d80260800184e08a8c13233ed84e6400b0321a05b556059ca929ba7a11ffbabcd31229a5835cfaf9aaf31138181ad9f0dd4ac235cb24fb56996bf94b0395fa14596f653a82e9ce783dcb4fe48ee1fba201546dfc6d904fee5418d2c90735d61189bb6e4b2b24d18dfff06c784e43f1c36c4b54c5100b9f09bbaced61d3f65fbc6b6ee478277e9a7321a59de9ebd8ce2fe94e60881162f74920bbf7f03997cf62d250a585dcf909b1a2754b53d935a31b48a28ac522ba273d7d90173d365d20fb16367b9a71526e337113fa585c23920aed8fb3f0078dea555f47418655230ed0e4087e7cf8b20883f8e34f1d58cfd0d461c05bcf4074391c79ae8bcaf6fb4e5ac270a69f7c98abb9fd3c2fbb989a39f8497e000b32ca377039c806766fe7eda55b67515599e485b8a0221d44322332bdee6753d8fa15180fd8d575aa702d290439176ce28e89f78f203df0087590d5672ba762bec02654103de24beec5590968d98f51759b7c3b0fd3374e7d090cbd7b8c25af1764e1b2ccdcfcc690c6209fccb8a206a88ec2e37cb351a89a836b54901254e727005dd6268da1e74c74e6d98a4beb34deea1372206a746f78ec2259e86e8f92dbaaaa748b5367da9955885a2c1bf1bec9fda5851ab9a0d3fbd529957b811b68dde1adac57acdf2ec0a41ac6ac187c7c1b712f8571fdcfbd62bc0e81814091fab4f41faf4ca136e507d24302b85e7f4d7d1cb233296dc45e9403a4de0838276a4d7b7ed8a3eafa106079ea21e2c1383ba3d14174f758eea8a19508d88b8d15f5ff2e6b2598d15c972c69aa61731efc382a942eaf0f6786ac1bfb916ce2bbd4cf53214cd54c71ba0c33047b17056b7dd2724810974b5bd13ae7df4d1240f61ff7ba4d1fdccfc457d4656ecd458486b6551a89a47711ea1a4c19da4ab49223359830083a7b1583c4a484f8b9a31273f46cca66ef3cd3402dc99e6220639991b7df8ea5a15a85fa5f9143bd65ded851f69dc47683cb007b552662586be2b1acd741ebc13d77635b07c9f98f459315a060ef1c97c1812ea69037ea72e2faaca0a61ec05ebc16600ffa856d7e0fac;
    localparam SPI_1 = 10000'h5e2b8ea5f31bfede8ea37db971d2af2fee2d0c0e7f508e4da88afeaf10d3a91efefd49857be3ba2c13c8c5d0b8f44c5542328adf5c8411e1ac3327bf87f233ecd1d2d18245797c0b664ee9adda0c01c7983ee095b36148cddb9abf2cb44e1909fc62917bd7e8f89f770fda92c6b44b96af632e4dc1baacd951ba31cfbb65a6eba9ab7d1c15c4dc2ad137b856a5805d7d2a009cde02744761f23a9ef3276f6cd0088cbb947167295080045c71d4ea7cc391d78078dfe0d2db9a179331da25515e7f99a0eafbd86f06ec0b48aa4f246c814a8fa862417297e403e9bfc213dd7bfe1cb749b39e4b8b65fc01da1a194f37591a239b508abfd4385cfce387644c3ce3234442902831cc7862adc9675ad9038a0a7d5ed055e50538d4c6f8e14015f1f053175b444d28533dcab899ab6d9109b11216a3dd7413b75a3d21d06d6463fb3e98fea9526ddafe79c0999b8ab456bbe52b3a8608babbf693a73e1f8a0320f1c93b2c4dc829e3c92f9fec03664b0095e012d947d0c5cf845ac314445c4034b06b245fb9d25c92ac4d951b050dcd86ce260544d724013287b5e09d52286a4997edff279195515eb977d30dcc4b8cfac32c0e0ebc4f8c9f686c963592a4679b82215e6883995d485a28210f85d19f9f42f40a4afd0fafb9ba690aa2910430d4aae5c47cbcafff3b0b93f4ab8504f68a8f94070e2dce7f8c668daa815f5b6e6c02544585871a28d249f884f872f2c31963abe50b526776eb2c8cf54f356321fd239d226b5e4ba15f919feab296348d94d83c9e68e9217f1bc7abd43bb67386cb1bb3beab6acb079f6150cc0c13e169357a2a8a0d5434b8a3f1241b53fd82db269bc17a6250bb5a588bcfbd13e4a8a76824adc55a23e992281254db9044f701962003b9c0d8c4f11e0b69be555f8bf585213ae9b7b1b57c9e98b071c21353e6911f454a16ded4023e1fc99602065777db8a8e644c959f6c73a0300157f2a0df54cc3766a3fc6d7f7f77564bf377cf58674840d4a47626058bf07588eb4a691971e76796ef255b61a20f483e683bd3e4056067cdb737ac734cf535b28cbe9f0d9fd2d55a98896f3b9daca14853134c772f4dcbdb6bb6e804d406316e07e78cf0edea4e51eb1f1b8e33c5dc9b18181d475511ac66b9bf7fc69c28a625abd7cf46c8d3ee7c6454708348410921011be2a9efbd6e0aad2d1d49fa5500dc7ddf7c186db72fed59789b5633778da36c9f734512617223d0598df38af6307233c6f012e52380c84f391964f335b7958188929fb0aa07a6ffccee1b7b7adbb68301cf78eb7d1d0683793376bcf9a47607cea231204608ee1a01c59b4696e208629ace3a98a45ad2449ee763ed4a505542e2ee9c294a54da11d5602816b8fdb47ed5260fd73bbc815d463aa1a9f9221808dcf7c5c3d7b33b73a70bff485432dcf01067b1b6389242f0a6ab77d7bca7c138c1f4e71c0f7a2ba7a838b7ec84489871c985391e2b06a65af6a712bccc39cfe8e9bd9b78f8025ada66fd98c7550743077e42101be12945986cac1d92813bfa5c614ce067e5fa6007c15bdc82a7363af98ebdc61acd073d0f52365c4a0641f0bd7ade8b893821c8a45cb4aa335e892ddb76afa2968998dd661faeccb7e8ecc3974955e85744de2ed3974af414cc560d8582777f16a64006ea1a3b36070efbf22f098e1b7a0fbba48d6f15bdca6da08aa8a481e4642b5b0004747f937a80204d68f92ad805fcaf2313fba26e3cfa3f811352f735433091a334;
    localparam SPI_2 = 10000'h7db6edf4152608c721810f45d8d8e8d95c4b3577b2bd855f326a3e39ed1235cc694efbd2227141b7397c2fd63758ec8f43705680c76ffc164a9238444ec0e2e8568e6bbc3eb50ef24661dc2a86d462e2fb98f753e1df933cdd41ea8c94a5bfddcc2e296345d49f747dfe5dd507c47b2844d850812cf7f54fb8c2ab2c458381f5236018f862338328eaabfe55807ad871a6f8e4120fe40aee1fad8ae1a3749f92fea088e071b81aa4089de21ac615be5ed5680977052d94a76e56a53f0bd0925bc0b94aa275af710987f1a3cc491c8f7f5edffa641d653bc3c6ac371ebcc2db8fe7bd1c223704ab75728829123945548e9bdac74f1f0ae36007b343b2f130809875ac272496136cdba60eb1910458cf2b793223f1c97149ea19612d1de9dafcce0c8539f896b85bd4d135182d7013e11745de864d97bfefae54d004c53c2fad331c3593e41aa6ce1e425e9017339ba9ba80a72ecca543ccf8a319550c149ec03f62ec8a72356a8d7efb47f8e728fac3e1b37fe5c77f62832667ccd807da0829d44efdc7929e033ac1c183313128d9ad09c2c5dd3f8af32a363ee39b09f05d9c5c522a91751b1092ef05c7c8f407bfc5671803ab362c840e7a1e7f6edd61227ab32abce24c715d6db3472f16729a32b4121bd8c8992e2f1beaf40e0b8dfd6abd02b5fe67f511f05de7736158edb1268d97edd1d0ce36d7b684d2fd27a0f8cf9954ec96ad5ab951c77967812604b3457bb525f3a86d54c9541193c301453feb2f7494fe9c7e7bf7c9a8c22bed19e4086d1d624a8bc0e2cc9b04981f2fc19c8c1f59480a35eb0a293e93f551d5588a5e47a30ec08082ad4e387cccf31fb044cdbe50fae85848c0b5f34d90fd3b5c2bde9b1b1a04774192aab20b158f9cc7413d2d775fcd70584f6ad73b96e4295dc8e56a7d4d5cee89c05c421d9ba4408c29f69b2110ac5008306a13d210007ae9ce7206826da54bc2969d67342ede7ed12f6df3eba0adc2bdac7f8df9b923ba1780758e1b66bd54dc6fed896e0c6ceffc3652ab1275a44efea2b97209b54525e4c22351715499e38fded34e844aee6bd972deca96e100bde6681973e038c0c66be931b02dfbcd0d7faa738451d376f2b9a5bcdb78306c8e4d5ed2742900e88e684b707eb439f5c1560873b972a4335fa3b655d2031661683c3e56f83496963fbc8f89cc8dab1f0969e385046968a6f6bd2eb76dad059497ff980bf0b52da386e51c9e9aebb18781acc5dce8c17858135387faaf287a346f025565364d908702b55e706d20a64bcb8d4330da25a6e911b877e52a4ad620a6c4c611b8afd4db0a1e40b84837b22fcb9fa07956659c13641ecb14fa93f406ae0409e62cd9efd656afeb157b941435b9cf310a628b63567e96a9793061b91a25497a881633096541b14b03df533e6fa3ddf77b50e309e115f147ead67d6c86768760eea817c0ec331d950ea3cc33b7fc51f777f36c89722e17ca8a4e1f8fabeadd5b50b0d55ef0c9496903ae176e530ac4b8f9f6a5699a8f0d2a65e3dc211d3592d4211e1bb619e5137ebdb1557dbc23dd006fe45da46038851741fab0ad1f839e28851323442a29b74dd4d28fce08c8f8000c64d083812eb6849ac042b047e51e7a70803527ec7ed822e74b2c0ad98a8c0a120aee11dcd93591c5e71eef08a9babbb32aebfc616a17a68657541b6ff169f5cae419c44ef380013e7c4b63d6cb71e8cc5f815813be04be0d96bc9159fa249a2cc3239533fb61b85aa16f0c5d;
    localparam SPI_3 = 10000'h742d7852e81f8202e702b528cdc916d4c4ba792d5fb44a1f721ec3ccf002f53da5da8eef3f610564c6a2be9e8bd7191e1c6e2fda729ca4d8648cac1b5745e265052d7839b889551391855380496b98b11f94c964f39b9282b04caa6d9730d49828a7068be28c8818715e0c9bf36ad733cd617a47e71c24f38febda4669fb621d1d971fe8062500f8f371bd101c2469bb8841c83407bd3804c01416ce77269b2192523fb6524aeca2815e539b12b6857c6fc236702c1b7f1d57a445f34c413899ffa60962cb36a91c8778fe71fb79e8b21ca2bb21e24b3fa7a53604b78129d53c51eb59804dd2a7d0265f31ea8d6b0d5f90e8cddc9bdff0025a7d889c8c323ab257179ee56d832741892a171d74d82fd49032f4909dfce15e69d44530df7fc91100f281856935ff310e5b505be57d420aca20a17c9bb55f59249668d24323cba0a3af2e74a586afa577fbc2b9ac2b32ecf8aea289aad673b7966ea079822179788db6382e35fd06b03be3e28faca026ca94b3f1db5fa0f2bd2ef9a07dfc9b550a276bdac2b7de05dc7bdee7ec32dac86d7944115f211b987157e89e4a95e3791b6600fe7620e05fcfa1598c130f66c51063c7472600751dcbc0566c8468a3198a5a23bde5a3590356f7bf3843fb5e9cb1e177dcc04babf472fecbcda2d28733e2ad8f1a1626cb36c0eba7cf04e5366cf02a40fbd07897daa1c7b26d9b052ce88303fa6eb322489cd2e2341c45288352e8f378c63f44fefd2815244da10b1738890375b1bb5de205c334fc1b922aa32f8030ed9ff9e5fad5f2238783ffe1f1a17a5f97086346c0da8ab5b6cfe5f13e4b6e9241c8afd882b3158fdd761d7773c46ca88d55c0456c8bfaceb0d782e503e2421b9f3df560b6b215356e8be950ce58f8de95d83a6339d56acfba25511ae67ee49876477042b8856ee1193ca9cf4eefecee044eb3e83095ee281a7e5d387b30749ef01e7ecc5403f221081d0724b0fda9ed220c2b46020cdd1d9fb5a05c59beb6b93a8ee14dbe8830d4491ac17643047a52303835b08be719102c76fe85bce8d61a2d02a638d29d9bb62d5f736b54743ca95e5346e4659d205c6f3e42f8dbbe07c667e266308c20fa771e8f88b117e5f8df51d6d2528c8ee739a546ca119e314cfbe75132569075196e3b4401d357404b93914a672273968706c9fe805f0dc2903054033f681435f3dae30666bfa55c669140dc4a07968f16e6e5bdcb17a7d98161c2ea54d63e63f0a82d4145383bdff07286447366518bf285265325a239a99a8ca38f50be71f50fe842e406a49d8e9e3817e81c552a24cb5a25159be39dc38bc3d232ef742a1bb05dd11ba930cc12fe56d0be34680a06ddff605c5e1b759b371835b3a2a8ac58183d5c93cab627b0aeb38f204a4b1dd2c5b30b82d64a27d88f5ca3dbdf15d522b9e9ca154e0dd163dfd75f7d3884cba0f2563d450ce6cde47678d416867c50c82ae628fb1add02c03ef577fffbf69d4c947b1d320dd286b23fa372f01d472428349b1a4dd1d7eeed086db699b013184d1f2f245562215260f6ea7842f46bb1595a126426496d7bf9d4db1ceeba7f9fdee9229a0f940c212eea187547a29169240ba84d3b89cd4caf54e9ee946d1d5ef1c73672d0e55e762ed78d1bc03fc698b7d53cdfc47b49d0222175d658ceb7eb7f8f8716c909a33c2a7eb0f9fc56655e3f25864d7a32b7dc72196dd89a526730fbbac58437b8fcfebe8ba4142e4aa5fdb2810b30693ce01805dc8cea;
    localparam SPI_4 = 10000'hd9d99dabfca7ddc341a101633da7c13367d57a3829e73fb8d11e294708d51135a2f0a30f5d14fcc1030dfd491c518ce5be563b81e47e04978aa5a2c6799cbe1509af930f745a2dcc04b91f820a140228a33ec56be68abea561e157ed33627e5b9562a45d1020023fd7ceb0886f65c1c86c167cd8e9ff55e340a007869185a664c755f0d6fac4a6f84161352530428e0d23c6b62382474326368c88519cc43dcb9b15e8be22af26b94ec99dfb5ca6aea96c207438bacd4f50cb1d5451ecef3a99dc50c26f2ba9c22ab0075d91d2b481d205801f2d97d8aa857f2c9790052d7fb8c1eea20fd4c10858e5b27dcb997eeab3d8c60c659b37602186de9823f620ea2a9589613b95966ad9dd8a7244b5f49a3218494bd18877ac88e0234929d76c115fb590e70275b03f09d378ca2e4d29ae436cadfc4905bf5f4d59af59bf06b7490ecdda6504e30371b4d364eadd491d9df4443f10e72dda8f25bf935c3e2bd1c63f3cd6b05e067078194503bbaed782bc50929c4df2adf53196cfd0a9da97738afbff12e47f4eec816822f70aeecef64283a123a2b7007b82a0a0c006989f55d4440d31aabe31ccb1090b819bd87b7e887a7cb7f069b277f1fdfa9525e7625cc6463cd8dc67574ee086361b1649ed864d2e46ea8f678561da746299ee6bc118706ca9f349bafae9bd52d0703382130e147d03d9034cd71a0ddad98769f032c39ddce3eb0d8d0abd733244463e40e9f2a39d05b43450ef3bea9cc9d8f23cb863b24a3a42323c610a5a59572d889c9679a380af9ce1f1481c2c8f1001739efd0bbc5ca541963d945a7d35699838d20311ad444f3bfbdbec8749048419d87c32328ff26197a6f72fb1c5af2e19629b0270223f9562758c70d04fcf29ab3ea8155319d589e671a54a0a8e4a826fbe79a68c908911284ac3727f15f6b190d9452a21e57a151a028ee3adda67088c13ec6ee847aa8850ccd3b410a30c38529aac6bb399c7cff219dead6779ce2513ffc2f9f757624ffda6a83fc3ec3db7e7a4d080d3445e992e3f7110ba6ea21d6a6d85f5fae6635ff74c756b0b722df36d5252cdb522ef2e1bb55559a943a9bedfdfd026d232ab874f9889539419a2a747c6d60cb0b5dfb5279beed73dca53381c8f7af28e2d932ba1f399a1ececf2df393960adddd57e6f89d5bf58c695db7f2c04a3d83598b218e98a43e149fceada0a1b9b94c0480a282a5504bd3e69c7f803fea37cb8e7d4511a3231b53570f0a33a1f26417a4b979b3f3dd9d51c09dc80aff90bc344db99ec715460d923f1e04fc95763db70b6611a8412d081318829ea408db7499bf9c2f8bd45e1ee195ff3cd83e8b5c15f1646fb9bfc917dd0b9e82449ed855dfbe9f497c57c37817b7da7aab52c8ba8b341f1516f6024701a81ed155b66513cb76983cd7717f183f3aa800e6a246fc00f0a745e19aeb56d955e6b931a50761dc5969ebed26c02c5f5b961e52d31c0540ad2abf7057ca051425a663d01fbf3eff4c8d57e37373702a785df9bc079b03947eac04995ba0c282916663ce4013eeeb4675b538fd0861ae666e27ae80e45785fa8061b48c5a96307d1a87b9694b148eb9d6e12805fbee4daf234b290f48c86f95ee797a453faecf67352aebf610375c2b5a02c58fed1ecbea3ba0636fc1626fe96306cd23d7809ec809db860973fdce038574ff036761a5799a690221594a9a890955dba8c835fe46c22974c06ea2a3a268ec18f28c66deea947f20258910f5b0ea2e6f9;
    localparam SPI_5 = 10000'h55f0bb97ab460a09015b03445fd329ee4648997514b4e9eb0963604ecfc679a3cfefbf2abbe8c8111866f8e370eb31d117e69559529d40ea6f78689fac736e9b60c6cd6b8b64f5150c9ecdae22ac5997c0d19276295beb272354b031acb89cf2ea0abd53b1190fd88ee492378602e9773045bd48f3ffbd0be619a1ee6f906d78c13d3ae90fd04201f9db3a3ad6220f7030e5692883eb0a374d4da8251fe5754204900a5ea78ea00741f5f0045a3cf52bfc6583baed895f17816cff4892b0223ebee445c410e9ce1905837d026e6338ef4943f194d94caabc222ec69a4751ec3b74bfb5233303b91896fd6ec29eb5fb66edc2c0442987876b558d5151dd78975072d11c16f6d57d3c5e907a0585d39eb2cde432851eaf307438d0becbccf2a8abcd858d93ba928ccbd86ca8fa800f4fdbd6f739046bfe2943f5dd80e04e78403c90cac1877434d6dd410a756a9df227c87416876085ced10d436752046a321fe9f3fd4fd6a3e6f5dcd1afa8d678ad6605c6d3499339b921d92f6e196c2efa9daf6481440c7b8229b860d64adfe57a56e370834bf7c833486a3e7ddc385589921ebef5ee21ab593e4c9555035b8d39d5d252e142b52658998fb891f79a137eef19517a6f578cfe33c64dcd6e448fca17eaac0cb73d98e744add53d1b55027c36aa386e9cc2b9bdb96dea8e379e1441a8aeee83a40a481d5c9eb698bd77ebf32267cc4884f7d80f8b5f0cbd072e4e0172fa5d9c6727ce97e88b6528d36e549ccb63dc64514317ec4eef572105bc50fb7be73b05abf81efcef7c79564faeb637b77eee87b609ada26f58ab524313e883086463951613e75354c0bfec8ddc0aac977a13a677ea8d30d2f41022393892f5dc16415f64d3717ec5f406494605851258cc0103a8e0d3c0d6e0fccd9258f58bb87520da3cc57eb9890222696cc0470daa4c5d32d5db6a5ac5c57d3248f30a5b1bbc30363610a4ed15ab6e23332dd9100dccedf7f804bcf9d43f1f50b1209e9a38ba113c7b659bf1748f215ba2eb270b06ae8e28ecd9afe9a04c11e1a5593bf5868de1b7b2cb923080434bd9f7c5ee96bdea129d9237a3c44253f1690651bb6e2274ceba567f79899e821fb42141fe149afd608f5187f72036c4e6cbe3ed3bb55c5fa2186587caa2a0f871b97de3718c076d9917170066e9fa58a98db2039d4924418fef0bfe5a6a4afb5c18558f7dd5a1d0ffee57b31590d6c33a7d8ce44a14be4534bd31b74b728433a1e2c38f72d03047a9619a122a2dc1db04e08d6422e293f94ccacbc8c34ead263d0917791bb49e8e540142dbfd1730eeabb910d8ade10fef0a052f21c3b130a9ed18a6e1ba9a3a6e81f6576488ad1e79ec9ef1308f5ceadad23581a8bb77b251122ecc4c4204a343bbbcd6dfb6e6a1e71d44aa4786f389840851ccd258484d231d2fdc3d0baa3a01877e19989b01984c746813af6314b76456ecc4eea94aee7e909ea470cc7c4d5fbd201db9876b7c7b29cecf8fd8e504a0e33ad0589ad8375b0be59916506bc587ef21a93d3d1ce15b0f13d86505f99c873619f75cc496aa25e553b1346c76c8b5f923a895d1a9af968cc9d0567031e299cbe27e80e202a288e78aa78879f257f02a0f7a72b9a660f40153178fd12d82f38a513cc263aa25154d35824281477525393e229cb20ea623b16a4a8d7b3cbc09142cbf7753d3d7b04d5282564ac997f1786d49dda56909fe96038b67cddae7b8c514a59b8d66506fbb0ae9c28344c9e01c96;

    localparam NUM_SPV = 64;
    localparam SPV_0 = 10000'hde3e35c39ff9941d9b59124b11e9ace6a9854343d3b0ac7a69581622e8e769430071e059cd1b03aa89e99163a479561bc6dc044a593a96bca97d319af6309eb406744f687f62daf4fdc46acf33b451b647f517478e2189ea1b2ec30b96c50ab694bc8a0c5cb679048ede91e77f7f816417d55ee33d0c002d66e98e9ad753c7b4d2064297d780a8810a3b64fdbe9e7fea46f2c813560144283e6d90b0bb364771cdbf8d31c8d809f68fc7a105e7c3bd18b73dd08c9f5ec821b1d9e731212f26905ee853edb7136ad6eda62facfa2ecdc76ffc1c89ecf8536f3fc7ccea5328036da1dd687d9e61bfd42f380e1385d5f18d5c50c23f2d1d5abdef0df9602752f8efabe8e1660209342abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_1 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcfff3b0ac7a69581622e8e769430071e059cd1b03aa89e99163a479561bc6dc044a593a96bca97d319af6309eb406744f687f62daf4fdc46acf33b451b647f517478e2189ea1b2ec30b96c50ab694bc8a0c5cb679048ede91e77f7f816417d55ee33d0c002d66e98e9ad753c7b4d2064297d780a8810a3b64fdbe9e7fea46f2c813560144283e6d90b0bb364771cdbf8d31c8d809f68fc7a105e7c3bd18b73dd08c9f5ec821b1d9e731212f26905ee853edb7136ad6eda62facfa2ecdc76ffc1c89ecf8536f3fc7ccea5328036da1dd687d9e61bfd42f380e1385d5f18d5c50c23f2d1d5abdef0df9602752f8efabe8e1660209342abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_2 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4c00000699163a479561bc6dc044a593a96bca97d319af6309eb406744f687f62daf4fdc46acf33b451b647f517478e2189ea1b2ec30b96c50ab694bc8a0c5cb679048ede91e77f7f816417d55ee33d0c002d66e98e9ad753c7b4d2064297d780a8810a3b64fdbe9e7fea46f2c813560144283e6d90b0bb364771cdbf8d31c8d809f68fc7a105e7c3bd18b73dd08c9f5ec821b1d9e731212f26905ee853edb7136ad6eda62facfa2ecdc76ffc1c89ecf8536f3fc7ccea5328036da1dd687d9e61bfd42f380e1385d5f18d5c50c23f2d1d5abdef0df9602752f8efabe8e1660209342abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_3 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435680000000309eb406744f687f62daf4fdc46acf33b451b647f517478e2189ea1b2ec30b96c50ab694bc8a0c5cb679048ede91e77f7f816417d55ee33d0c002d66e98e9ad753c7b4d2064297d780a8810a3b64fdbe9e7fea46f2c813560144283e6d90b0bb364771cdbf8d31c8d809f68fc7a105e7c3bd18b73dd08c9f5ec821b1d9e731212f26905ee853edb7136ad6eda62facfa2ecdc76ffc1c89ecf8536f3fc7ccea5328036da1dd687d9e61bfd42f380e1385d5f18d5c50c23f2d1d5abdef0df9602752f8efabe8e1660209342abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_4 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bac0647f517478e2189ea1b2ec30b96c50ab694bc8a0c5cb679048ede91e77f7f816417d55ee33d0c002d66e98e9ad753c7b4d2064297d780a8810a3b64fdbe9e7fea46f2c813560144283e6d90b0bb364771cdbf8d31c8d809f68fc7a105e7c3bd18b73dd08c9f5ec821b1d9e731212f26905ee853edb7136ad6eda62facfa2ecdc76ffc1c89ecf8536f3fc7ccea5328036da1dd687d9e61bfd42f380e1385d5f18d5c50c23f2d1d5abdef0df9602752f8efabe8e1660209342abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_5 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4340000cb679048ede91e77f7f816417d55ee33d0c002d66e98e9ad753c7b4d2064297d780a8810a3b64fdbe9e7fea46f2c813560144283e6d90b0bb364771cdbf8d31c8d809f68fc7a105e7c3bd18b73dd08c9f5ec821b1d9e731212f26905ee853edb7136ad6eda62facfa2ecdc76ffc1c89ecf8536f3fc7ccea5328036da1dd687d9e61bfd42f380e1385d5f18d5c50c23f2d1d5abdef0df9602752f8efabe8e1660209342abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_6 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3f80166e98e9ad753c7b4d2064297d780a8810a3b64fdbe9e7fea46f2c813560144283e6d90b0bb364771cdbf8d31c8d809f68fc7a105e7c3bd18b73dd08c9f5ec821b1d9e731212f26905ee853edb7136ad6eda62facfa2ecdc76ffc1c89ecf8536f3fc7ccea5328036da1dd687d9e61bfd42f380e1385d5f18d5c50c23f2d1d5abdef0df9602752f8efabe8e1660209342abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_7 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef4000000be9e7fea46f2c813560144283e6d90b0bb364771cdbf8d31c8d809f68fc7a105e7c3bd18b73dd08c9f5ec821b1d9e731212f26905ee853edb7136ad6eda62facfa2ecdc76ffc1c89ecf8536f3fc7ccea5328036da1dd687d9e61bfd42f380e1385d5f18d5c50c23f2d1d5abdef0df9602752f8efabe8e1660209342abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_8 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44000000cdbf8d31c8d809f68fc7a105e7c3bd18b73dd08c9f5ec821b1d9e731212f26905ee853edb7136ad6eda62facfa2ecdc76ffc1c89ecf8536f3fc7ccea5328036da1dd687d9e61bfd42f380e1385d5f18d5c50c23f2d1d5abdef0df9602752f8efabe8e1660209342abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_9 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c2388c9f5ec821b1d9e731212f26905ee853edb7136ad6eda62facfa2ecdc76ffc1c89ecf8536f3fc7ccea5328036da1dd687d9e61bfd42f380e1385d5f18d5c50c23f2d1d5abdef0df9602752f8efabe8e1660209342abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_10 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ecaad6eda62facfa2ecdc76ffc1c89ecf8536f3fc7ccea5328036da1dd687d9e61bfd42f380e1385d5f18d5c50c23f2d1d5abdef0df9602752f8efabe8e1660209342abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_11 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307acbfffffffffffff836da1dd687d9e61bfd42f380e1385d5f18d5c50c23f2d1d5abdef0df9602752f8efabe8e1660209342abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_12 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd1ffffffffffffffffffe23f2d1d5abdef0df9602752f8efabe8e1660209342abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_13 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fdffffffffffffffffffffe2abe3f546f9062a4171c1ac3e2850d7697f93d9af3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_14 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3fffffffffffffffffffff3daafb231cbae6d5485eb7a65d284b03a993f3b6322be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_15 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345197fffffffffffffffffffffffffff2be3445b39da7992f66110cfbcfe2477f059e019de4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_16 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c62fffffffffffffffffffffffffffffff4eef62d2f56f3a098e5ed197f436b0bcfdbb6b563690f5c0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_17 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109dffffffffffffffffffffffffffffffffffffffffe0d10b906b531271ed06de29efc53c832abb8b232df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_18 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9ffffffffffffffffffffffffffffffffffffffffffffe32df3c2e1ef01cb9b16b67f745605278fde3d9369f84d1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_19 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54fffffffffffffffffffffffffffffffffffffffffffffffcd1249a41a96422a0a344c27842acbb103d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_20 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad8707fffffffffffffffffffffffffffffffffffffffffe3d49e0c3c0579c6604598cccf4efb9aea6871d5a2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_21 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2bffffffffffffffffffffffffffffffffffffa2bc4ade9075568a0ca3a01984d7996be9771ac0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_22 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43ffffffffffffffffffffffffffffffffffe0d2e95cdf20440acdfff02b66e419314bae2ae28aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_23 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a7fffffffffffffffffffffffffffffffa8aab3e065e811be241a2cb13d3726eed674362b244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_24 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9fffffffffffffffffffffffffffffeb244649449308e0e13c0e599e07805dc4dcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_25 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71fffffffffffffffffffdcac79e443852f2b67eaf4a531cb346f29ab32be772801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_26 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150ffffffffffffffffffffff801be869c034b51534ad4ac05c9f4efe051427d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_27 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb53fffffffffffffffe27d0b224657bd41d91f09fd4bd5c31dd2412700f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_28 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b7fffffffffffff8f3d6ab5b51b8e06b2b0fff1102b83a68b9b44680eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_29 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eeffffffffffffffe0eca1ba0d330e787d9a86b6fd9697591113cf5060a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_30 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026fffffffffffff60a4b083512e71c10163a6544a4fa52f34dd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_31 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cffd06b2dffb9a5b8588178b7bb5bb8690f646a63d32337c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_32 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09bbfffffffb7c4be493edc3ec8a3fbbcfe380e90e03da607c6fc297e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_33 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f17ffffffffffffffd7e23a3a1370c382d759681f37404fb9f3b655f47787dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_34 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8ffffffffffffffffc7dde561d6e3055bf1de7defe6f80c79f9f3b70a148e20e32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_35 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e3ffffffffffffffffffffffffffee32fe7421c4de2c1d5c2efde50aecc1e2d6465e3b75f040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_36 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bdefffffffffffffffffffffffffffffffffdf040fa2d90c1423adc493856660ab04258751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_37 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf7ffffffffffffffffffffffffffff8751172a58f174a4f9d9c71db640f061287cae89c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_38 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b3fffffffffffffffffffffc9c324f86557df323a0f211295579d32d16f049612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_39 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5fffffffffffffffffffff612ae0b23dd9e8413fdd801f64c87f06e5061c620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_40 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec022fffffffffffffffffe620b836608f89e90c39a2498f81f365d5e354ce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_41 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e1ffffffffcce0b2472cf15dd569c9274ef77a5ccb1ca9b7e44412892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_42 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885bfffffffffffff92892ab3b5e4e489220346310a2371807fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_43 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8fb94b03e485bdca6955d25c8b578a36d3366e5aa9c3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_44 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991affff3f4527d8c4ff11d2e705b2bf6d5ae08b95dd24561c309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_45 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746ffffffffe309eb64e7c992cf8792300121c21b40a5c0d26b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_46 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a30006b789e98e4d055b598086dde765a781dd66a79f7dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_47 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e229958477dc22fe6b70be5ef98835fd57ac1661a6f4adc050b6d158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_48 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e593ffffffffed158c19b7797b2c599729105e1d7294592bf608159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_49 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6bbffffffc159f6337086a1ed979c5a19a0d8684020abf7956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_50 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf5407956eeeee3d3dcf485bef2ed83c549d36bd6a3e4c4e5b04961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_51 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf54086a911111c2c230b7a410d127c3ab62c97ffffffffffff4961c4547690f1ab4642af7c1a7dc6156b95d6cc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_52 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf54086a911111c2c230b7a410d127c3ab62c94295c1b3b1a4fb69e3bab896f0e54b9bd5083e583fffffffffffc7382ebfb9ca761983187a23ba58e9788a470800df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_53 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf54086a911111c2c230b7a410d127c3ab62c94295c1b3b1a4fb69e3bab896f0e54b9bd5083e58239ea946a29338c7d140463589e67ce785dc45afffffffffffc0df12ca0e5f43e1c6d036c61e42872e677a8127fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_54 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf54086a911111c2c230b7a410d127c3ab62c94295c1b3b1a4fb69e3bab896f0e54b9bd5083e58239ea946a29338c7d140463589e67ce785dc45a7168775b8f7ff20ed35f1a0bc1e392fc939e1bd78d19bfffd27fd4c643438e4202dc2c9f551097d926f7b83870ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_55 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf54086a911111c2c230b7a410d127c3ab62c94295c1b3b1a4fb69e3bab896f0e54b9bd5083e58239ea946a29338c7d140463589e67ce785dc45a7168775b8f7ff20ed35f1a0bc1e392fc939e1bd78d198857ed802b39bcbc71bdfd23d360aaef6826d9084ffc70ad1b2040365d6eaafe4622b4f1f6f2e64c9b0668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_56 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf54086a911111c2c230b7a410d127c3ab62c94295c1b3b1a4fb69e3bab896f0e54b9bd5083e58239ea946a29338c7d140463589e67ce785dc45a7168775b8f7ff20ed35f1a0bc1e392fc939e1bd78d198857ed802b39bcbc71bdfd23d360aaef6826d90847c78f52e4dfbfc9a2915501b9dd4b0e090d19b367c668cbd7eb161ae4ed5797ac2c5527329f28949079aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_57 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf54086a911111c2c230b7a410d127c3ab62c94295c1b3b1a4fb69e3bab896f0e54b9bd5083e58239ea946a29338c7d140463589e67ce785dc45a7168775b8f7ff20ed35f1a0bc1e392fc939e1bd78d198857ed802b39bcbc71bdfd23d360aaef6826d90847c78f52e4dfbfc9a2915501b9dd4b0e090d19b364f997342814e9e51b12a86853d3aad8cd60d76bff79aab654732fc6cedfaeba8c5c247c0f4084d844faa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_58 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf54086a911111c2c230b7a410d127c3ab62c94295c1b3b1a4fb69e3bab896f0e54b9bd5083e58239ea946a29338c7d140463589e67ce785dc45a7168775b8f7ff20ed35f1a0bc1e392fc939e1bd78d198857ed802b39bcbc71bdfd23d360aaef6826d90847c78f52e4dfbfc9a2915501b9dd4b0e090d19b364f997342814e9e51b12a86853d3aad8cd60d76b6f865549ab8cd0393120514573a3db83f0bf7b27fffaa01d406e946c26fc8e9cdda2072cebe633c54df08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_59 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf54086a911111c2c230b7a410d127c3ab62c94295c1b3b1a4fb69e3bab896f0e54b9bd5083e58239ea946a29338c7d140463589e67ce785dc45a7168775b8f7ff20ed35f1a0bc1e392fc939e1bd78d198857ed802b39bcbc71bdfd23d360aaef6826d90847c78f52e4dfbfc9a2915501b9dd4b0e090d19b364f997342814e9e51b12a86853d3aad8cd60d76b6f865549ab8cd0393120514573a3db83f0bf7b27bb055fe2bf916b93d9037163225df8d31419cc3abdf08739a08f5e9efc149ecbec983c7ac3b4f87920420990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_60 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf54086a911111c2c230b7a410d127c3ab62c94295c1b3b1a4fb69e3bab896f0e54b9bd5083e58239ea946a29338c7d140463589e67ce785dc45a7168775b8f7ff20ed35f1a0bc1e392fc939e1bd78d198857ed802b39bcbc71bdfd23d360aaef6826d90847c78f52e4dfbfc9a2915501b9dd4b0e090d19b364f997342814e9e51b12a86853d3aad8cd60d76b6f865549ab8cd0393120514573a3db83f0bf7b27bb055fe2bf916b93d9037163225df8d31419cc3ab20f78c65f70a16103eb61341367c3853c4b0fffffc20990517b1ffed2512add6cb192cb558ce4c81cc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_61 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf54086a911111c2c230b7a410d127c3ab62c94295c1b3b1a4fb69e3bab896f0e54b9bd5083e58239ea946a29338c7d140463589e67ce785dc45a7168775b8f7ff20ed35f1a0bc1e392fc939e1bd78d198857ed802b39bcbc71bdfd23d360aaef6826d90847c78f52e4dfbfc9a2915501b9dd4b0e090d19b364f997342814e9e51b12a86853d3aad8cd60d76b6f865549ab8cd0393120514573a3db83f0bf7b27bb055fe2bf916b93d9037163225df8d31419cc3ab20f78c65f70a16103eb61341367c3853c4b0786dfbdf66fae84e0012daed522934e6d34aa731b37dcc7a9d96cf24868b2c296a1a5b887a7a5b6a4b1acdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_62 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf54086a911111c2c230b7a410d127c3ab62c94295c1b3b1a4fb69e3bab896f0e54b9bd5083e58239ea946a29338c7d140463589e67ce785dc45a7168775b8f7ff20ed35f1a0bc1e392fc939e1bd78d198857ed802b39bcbc71bdfd23d360aaef6826d90847c78f52e4dfbfc9a2915501b9dd4b0e090d19b364f997342814e9e51b12a86853d3aad8cd60d76b6f865549ab8cd0393120514573a3db83f0bf7b27bb055fe2bf916b93d9037163225df8d31419cc3ab20f78c65f70a16103eb61341367c3853c4b0786dfbdf66fae84e0012daed522934e6d34aa731b37e3385626930db7974d3d695e5a4778585a495b4c2cdc92d719a595e449f20932d92eb4f891cf6d52;
    localparam SPV_63 = 10000'h21c1ca3c60066be264a6edb4ee165319567abcbc2c4f538596a7e9dd171896bcff8e1fa632e4fc5576166e9c5b86a9e43923fbb5a6c569435682ce6509cf614bf98bb097809d250b023b9530cc4bae49b80ae8b871de7615e4d13cf4693af5496b4375f3a34986fb71216e1880807e9be82aa11cc2f3ffd29916716528ac384b2df9bd68287f577ef5c49b0241618015b90d37eca9febbd7c1926f4f44c9b88e324072ce3727f60970385efa183c42e748c22f7360a137de4e2618ceded0d96fa117ac1248ec95291259d05305d132389003e3761307ac90c0383315acd7fc925e229782619e402bd0c7f1ec7a2a0e72a3af3dc0d2e2a54210f2069fd8ad071054171e99fdf6cbd541c0ab906f9d5be8e3e53c1d7af2896806c2650c25504dce345192ab7a14859a2d7b4fc566c0c49cdd41cbba4c625866d099eef304301db880fa61fe621b1109d2d0a90c5f671a12e680bc94f43024494a9c96f0a3f2ef46f94aced8e12f921d6103ac37cd54474dcd20c3d1e10fe3464e949808ba9fad87021c26c9607b2edb65be569bdd5f5cbb3d87bd5344efc2b61f3c3fa86399fba673330b1046515978e2a5d43b5216f8aa975f35c5fe67b2866941688e53f2d16a320dfbbf532000fd4991be6ceb451d51d7554c1f9a17ee41dbe5d34ec2c8d911298bc9d4dbb9b6bb6cf71f1ec3f1a661f87fa23b2353861bbc7ad0d498150b5ace34cb90d654cd4188d7fe417963fcb4aeacb52b53fa360b101faebd82f4ddb9a842be26e0f602b42a3ce22dbed8ff0c2954a4ae471f94d4f000eefd47c597464bb97f135e45f2ccf18782657949026968a6eeec30af9f5b4f7caed18e3efe9c59abb5b05ad0cb22f94d200465a47a77e874844a44796f09b959c2cdcc83b41b6c123c1375c044301c7f16f1fc259f83903d681dc5c5ec8f3c7d28a697e0c8bfb0460c49aa0b8878221a9e291cfaa40e2182101907f386060c48f5eb71df1cd018bde3b21d3e2a3d1021af5133e1d29b9a1c48a0fbf05d26f3ebdc523b6c7a999f54fbda78aee8d5a70e8b5b062638e249bf0f9ed78351763cdb079aa820cdc5f0deed6aa862cd2e90fb69ed51f4dc22617bec0227fe09b3780f91af9e39df47c99f707616f3c65db6707e0c9a2a1cab31f4db8d30ea22a9636d8b10885a334e356481bbbed76d54c4a1b1b76ddfcb9cef5dc8e7f8046b4fc1b7a423596aa2da374a875c92cc991a5563c0bad8273b00ee2d18fa4d4092a51f746a22dba9e3cf6149b18366d30786dcffede3de4bf5a3f2d948761671b2faa4a67f7922189a587e22995860823dd01948f41a10677ca02a853e99e590b523faf492ea73e6488684d3a668d6efa1e28d6ba6d409f7ea609cc8f795e126863a5e65f2797bfdf54086a911111c2c230b7a410d127c3ab62c94295c1b3b1a4fb69e3bab896f0e54b9bd5083e58239ea946a29338c7d140463589e67ce785dc45a7168775b8f7ff20ed35f1a0bc1e392fc939e1bd78d198857ed802b39bcbc71bdfd23d360aaef6826d90847c78f52e4dfbfc9a2915501b9dd4b0e090d19b364f997342814e9e51b12a86853d3aad8cd60d76b6f865549ab8cd0393120514573a3db83f0bf7b27bb055fe2bf916b93d9037163225df8d31419cc3ab20f78c65f70a16103eb61341367c3853c4b0786dfbdf66fae84e0012daed522934e6d34aa731b37e3385626930db7974d3d695e5a4778585a495b4e53236d28e65a6a1bb60df6cd26d14b076e3092ad;


    input [$clog2(NUM_CHS) - 1: 0] c;
    input [$clog2(NUM_SPI) - 1: 0] spi;
    input [$clog2(NUM_SPV) - 1: 0] spv;
    output logic [DIMENSIONS - 1:0] ch_hv;
    output logic [DIMENSIONS - 1:0] spi_hv;
    output logic [DIMENSIONS - 1:0] spv_hv;



    wire [NUM_CHS - 1: 0][DIMENSIONS - 1:0] ch_mem;
    wire [NUM_SPI - 1: 0][DIMENSIONS - 1:0] spi_mem;
    wire [NUM_SPV - 1: 0][DIMENSIONS - 1:0] spv_mem;


    assign ch_mem[0] = CH_0;
    assign ch_mem[1] = CH_1;
    assign ch_mem[2] = CH_2;
    assign ch_mem[3] = CH_3;
    assign ch_mem[4] = CH_4;
    assign ch_mem[5] = CH_5;
    assign ch_mem[6] = CH_6;
    assign ch_mem[7] = CH_7;
    assign ch_mem[8] = CH_8;
    assign ch_mem[9] = CH_9;
    assign ch_mem[10] = CH_10;
    assign ch_mem[11] = CH_11;
    assign ch_mem[12] = CH_12;
    assign ch_mem[13] = CH_13;
    assign ch_mem[14] = CH_14;
    assign ch_mem[15] = CH_15;
    assign ch_mem[16] = CH_16;

    assign spi_mem[0] = SPI_0;
    assign spi_mem[1] = SPI_1;
    assign spi_mem[2] = SPI_2;
    assign spi_mem[3] = SPI_3;
    assign spi_mem[4] = SPI_4;
    assign spi_mem[5] = SPI_5;

    assign spv_mem[0] = SPV_0;
    assign spv_mem[1] = SPV_1;
    assign spv_mem[2] = SPV_2;
    assign spv_mem[3] = SPV_3;
    assign spv_mem[4] = SPV_4;
    assign spv_mem[5] = SPV_5;
    assign spv_mem[6] = SPV_6;
    assign spv_mem[7] = SPV_7;
    assign spv_mem[8] = SPV_8;
    assign spv_mem[9] = SPV_9;
    assign spv_mem[10] = SPV_10;
    assign spv_mem[11] = SPV_11;
    assign spv_mem[12] = SPV_12;
    assign spv_mem[13] = SPV_13;
    assign spv_mem[14] = SPV_14;
    assign spv_mem[15] = SPV_15;
    assign spv_mem[16] = SPV_16;
    assign spv_mem[17] = SPV_17;
    assign spv_mem[18] = SPV_18;
    assign spv_mem[19] = SPV_19;
    assign spv_mem[20] = SPV_20;
    assign spv_mem[21] = SPV_21;
    assign spv_mem[22] = SPV_22;
    assign spv_mem[23] = SPV_23;
    assign spv_mem[24] = SPV_24;
    assign spv_mem[25] = SPV_25;
    assign spv_mem[26] = SPV_26;
    assign spv_mem[27] = SPV_27;
    assign spv_mem[28] = SPV_28;
    assign spv_mem[29] = SPV_29;
    assign spv_mem[30] = SPV_30;
    assign spv_mem[31] = SPV_31;
    assign spv_mem[32] = SPV_32;
    assign spv_mem[33] = SPV_33;
    assign spv_mem[34] = SPV_34;
    assign spv_mem[35] = SPV_35;
    assign spv_mem[36] = SPV_36;
    assign spv_mem[37] = SPV_37;
    assign spv_mem[38] = SPV_38;
    assign spv_mem[39] = SPV_39;
    assign spv_mem[40] = SPV_40;
    assign spv_mem[41] = SPV_41;
    assign spv_mem[42] = SPV_42;
    assign spv_mem[43] = SPV_43;
    assign spv_mem[44] = SPV_44;
    assign spv_mem[45] = SPV_45;
    assign spv_mem[46] = SPV_46;
    assign spv_mem[47] = SPV_47;
    assign spv_mem[48] = SPV_48;
    assign spv_mem[49] = SPV_49;
    assign spv_mem[50] = SPV_50;
    assign spv_mem[51] = SPV_51;
    assign spv_mem[52] = SPV_52;
    assign spv_mem[53] = SPV_53;
    assign spv_mem[54] = SPV_54;
    assign spv_mem[55] = SPV_55;
    assign spv_mem[56] = SPV_56;
    assign spv_mem[57] = SPV_57;
    assign spv_mem[58] = SPV_58;
    assign spv_mem[59] = SPV_59;
    assign spv_mem[60] = SPV_60;
    assign spv_mem[61] = SPV_61;
    assign spv_mem[62] = SPV_62;
    assign spv_mem[63] = SPV_63;

    always_comb begin
        ch_hv = ch_mem[c];
        spv_hv = spv_mem[spv];
        spi_hv = spi_mem[spi];
    end

endmodule