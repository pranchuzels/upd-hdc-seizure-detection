`timescale 1ns / 1ps
 
module tb_similarity_hf_mapped;
    localparam T = 10;  // clock period in ms

  // General Params
  localparam DIMENSIONS = 10000;

  // Port declarations
  reg clk;
  reg nrst;
  reg en;
  reg [DIMENSIONS - 1 : 0] hv;
  reg [DIMENSIONS - 1 : 0] ns_hv;
  reg [DIMENSIONS - 1 : 0] s_hv;
  wire out;
  wire label_out;

 
  similarity_hf #(
    .DIMENSIONS(DIMENSIONS)
  ) 
  u_similarity_hf(
        .clk(clk),
        .nrst(nrst),
        .en(en),
        .hv(hv),
        .ns_hv(ns_hv),
        .s_hv(s_hv),
        .out(out),
        .label_out(label_out)
    );

    // Clock
    always begin
        clk = 1'b1;
        #(T / 2);
        clk = 1'b0;
        #(T / 2);
    end

    initial begin
        // $vcdplusfile("tb_similarity.vpd");
        // $vcdpluson;
        $sdf_annotate("../mapped/similarity_hf_mapped.sdf", u_similarity_hf);
        nrst = 0;
        en = 0;
        hv = 0;
        ns_hv = 0;
        s_hv = 0;
        s_hv = ~s_hv;
        # (50000000 - 5)
        nrst = 1;
        en = 1;
        hv = 5'b00001;
        # (5 + 5)
        en = 0;
        # (50000000 - 5 - 5)
        en = 1;
        hv = 10000'hceec8d666e2132e1c2a669e8012a05ee5a74e15c0833feedd32b9ce714002c06914b6014e155f7927f0fdc9f38354d460f4ecc00b51691d434a00ebe8e5484123bf7d3347277c9052227be0ee96e351ae5a287e605224aca787e129a77e32b628d77f9bffb16f478660a3904a2a14c80cc6a8ac0c17fd12840db0a1e09ee8f83c315bf78ddcf312079a32fb9a181dba69b8a660b2df8fc976770564a1d2bd7645d3d68a953cd95ca50720ae0678f5e1459ae103ec6c018947dea42cd98301a48b2220390e761d57d7406c860d1e4c69e48d857d92f259791e8ae2cba0de6fdd1e5aac08462476a986a1b5643a904bb0079a48d562b5a75cef02cd4a5a50d87bd2e1031490f4af6c36f67f4b458c0f3f77116ca5ad0a6854c97b46dd4bf884c2c29dd39cf8749383cd783128108eadd1e5888ecd53b30336b871cfbc3c008492a40502a3e24627adb4d9c451d02ce6c57b237e6020fe94d4c73d9383068e7b67fb5fd54d57692f1f4c59d417732958fc38189617e065c6dadfe2a3a974088d6f00ee0efa9d3f83061e7488d1ff33d8b2207f3762b16e900adbae25583abd52750453163e802dd0d9586743f1688e3f6a0d9864dc54751747f00c3dba3aa5700123836f643d169e412e56f19a725b8a797cf8165c5bb623df7f30ab1787a11993bc3939898a83003835eacf8b13f45f7f0ff6702da5c20b76a5ff32706e9db982df03a9657a614188d8e34826fa5c131bd572fcb0ea0db42a0d271225112430b284e3da3a4e9858f2e40accb180591bf63eb62c807ef3a417897bbb6526de3ab0ecebb8a5ea97d5f779a8da2c135d5d6bf77d2881f9faf003cc6234de09f71935a1caef8a1972e10eeff54f4588fc5241cb65b915339c6acefdf5653195900e677e69c40075c8ceabca77c36a9b44dd5a078da855377c5aeaeb9513a6faa90cddde2d9c3adbe90cc710cbc2b699a4bab6d50298ffc3638bb23fdeaa95495bb882f4c241564fc2fcb23477896efb1ded875635f893cbc4e2b7138fc24bf3e464bd38b3ad8ec4be0afa6a85a1b988b3240aae0f49269fd5331b1b4681eb11a558a70bb9880078d14c88ffb900b2553a989f54e49b87b81d8a3ad58847d87f7a9f5286908bf7c29c80cdde546f17bb2fcee21a845dd91ba9f7c31e2a8e71872e532a57f41c2ecfe0fee20e6e8d314bd68d27870d47d1352811ec499cc0b24300411f442565273625fe26e11af3e67852b574863bed650c003e98560648db70dcc2b0f30ac5b9684f50e1c3265dfa11697ae827ebf114a2837c3021bf0294093090f2881d44a4c0105e9a48d3c0e0d08cbabfde3ec6a46b9bce69c2977a33335091685188252afe678c2c81c75ad6ed8700c49d5815dfb36e950d9ec0979287149c8a01abb86a20dd2645ba91d1239ccfa0850889d313218a247eee01adf0bba7f13d71f3ea4a5a0e7b3c076f17166362d82291f8081249606517d29c5ea52b27ac4612b59637752fe1da480d96e43645eda8b2ba50aa3b19a343a8765a936f0798e00cf0f234d285a16e662facf4110fffb40e32cbb1c468a404e925072592cf77ea8fc917d7245686b9a76919852f8379ed6d505a1f42b13ae49160e2b71d6dd88ce805c927c196c50df8f4ce5a2e70e7565c6555b226447c6491fb6220f6ceaaeabf51086fcfa0259ce63392fd682e402dcc8738378bb201b1bb4c0ee603a8cbd6634ff9b162bc882d136080745abf6f8d85afa54f875d18a3fca376abd10b31247a5f0;
        # (5 + 5)
        en = 0;
        # (50000000 - 5 - 5)
        en = 1;
        hv = 10000'hdfc8f6f8880169970491d765c95443cf702b5e153781cdd7f3e0f67c5f00a0b7b6bab8b4f718469b964da695efa99e663ef2b83246afe9d0d0b4175c17b4af8884461b14091834d45da579714223ed2a94c5fc7cfb28aa2d267865ce7c8701f7586c37c4db9e21b89bf4b3466e7cef079202f6bccabe3e390eb82cae4f704b1d4cac65005bdba199ac03a4c27f5d5fa2e3e94eb3746a36004440bed59150db6ad3f03f8fbcdd94af5ab861e0ec75c5844df2ba3e79a2851cacb553a25641bf45b43d41c0984c0fbf583fcf6a04b4a359a53a62de684d5dd7845809cdd5c6fa4934034f63e4128f411710b7792486e53af4717be3a4ca18bec514781965a54436cf1e4e82c2a4b72fbdcc08ede19c59a786867e573b9a9e385ef3f16da92d0f5d374f6ff1fe591db413aadec612b5d4e2c6224fc4399845bb47be65e63f7240a557ca064c1efc7f345aced097eb27e9a105f1eff8fc154e3974d401d6d492131e37a74cf8e950886339f9708cb477cc9d2954b5338fdc23055a0a543a7e8090bebd37182b3d1675057ac6e36efed229f4ffb5f152fb1980f8db011bd7e2498f8c960f69f9fd24172fc66002004bcb29c4fb5b1d8915db8a9d3e6c483f1277af9abf0b2d1a2384a85f484d7af609a88ea036dc3022269e07e08360ae9874426be499bf17b8f43e8617b1eec83e9ab32038a45242dacb6b25e52cd865df1ef0df30d4a6771e5b21c8d325ab6691e0d34df566a76597fcaf91d121622ffe06bb21458e751ef94e05e79feb354252c8f1565b4ffbe21d7353a155abaf1fe051b616381b628c96b6f6fab46470918d2e50bfad492c3a5761f08eb6f0c43519ac06d0c7a93b1d4cf579942938f919458cfed15f10134b8395c701a0db72b858219b698eb45ec30a9af379f2dff902617a02d8cfd3a0ed496520d293b537c24a305b68be6463746c2a5fec0b25e76e95162dab61dbc0b002e64a8b9d8ea03fa7f27f2d5a70ba18acb16abfbcdcc9a52182de16a8a89a0e7a84ca6096320fd816149ef0257a2c95dd2f2688b6951a0adae278544eacc42999144b2bbe44592e8643b8cd11f80ad68a89e6eb31baa8a5b604d691eb06895d14e85099df8e0928f70c1b5c420f8fb2223393884e571acc0bea85a090fb2bebb367889ed9c2d7dcfc19a8adb4f19f680a3d010b5d1fab7d2f9a88998287e5c8c9f4ac66615b55fb60d608dc6d55aab52ce4e48d8720168274354e39f121fb118d7f3bd84f53b7cfb581c5c7975ee20fab9ab5ade35d37e7ea6d7f8eb5c5662c80b5d5d5786ba55b56dd1fdc32404c7e1a6f0d656479ed15a617419a1f30ea6e241f4ff34c6bfaab408fe698b2c950399c3fbe4a0c9974c463af52e0efd70ff96ab456532a6e48d7af1cb2e50e0cc7e2aa0b055a892d659980991108bd661aa9ebd340638c61d9343cfa12448bc884beec62e85faef2e37279259d1dd994286f6cbfb2a1a89152066e52cd30276613dabafa6b195fdbac50b2c52fcb5a5ab1d2bd10b5a88f80f2727d4b1e47e8f3995d1df0a26f2b5746791193c1ab32e85f3d96824acbeadf6f1bd5754742366c6915c9742c3f1e572047ec1ec5ddcdc4124b4a8b6aec006aeb9cc8abab0a00653fd7f9f3a318f8c998f002314cd1b075717bdabef90b34a571650a8a3f71e003248e9e060f67c5a51847098ec4f4dc6046acfd5ce1860250cb37432c936af4385eeab03b18bc0c0b9801993ff71b33326d4f84ec0468919627721798d3b84319f6;
        # (5 + 5)
        en = 0;
        # (50000000 - 5 - 5)
        en = 1;
        hv = 0;
        hv = ~hv;
        # (5 + 5)
        en = 0;
        # (50000000 - 5)
        $finish;
    end
endmodule