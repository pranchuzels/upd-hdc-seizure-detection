`timescale 1ns / 1ps
module item_mem_1 ( // LBP
    c,
    l,
    ch_hv,
    lbp_hv
    
);
    // General params
    localparam DIMENSIONS = 10000;

    // Channel params
    localparam NUM_CHS = 17;
    localparam CH_0 = 10000'h385ece781dc2bccbd165b943df9f6c66b342c66c2874ae514e0711f121c41f048801feea276873b287bd12f502941a94be1d5f096e25de5e8302869cf77bcd54cfd2d567c57009926b1e29ed122d3749a60ab4bacd37df3243211580480e608ec4e592429b0d1813ab99ea6aaf8c41c9d8ea9896e3baa370797ae8d60df7548c8efd8b349e70a8f730fdd5dbcd3ad80b195b0f7f19e49b9b6f3e20e47646a8e58fe927df1657183795426abe022894cdb1daea13b3b99845b8afb3e1f1407726da678ac5c0ad293ae4e05310e3ac2644596229882bf2a82c245403f0455dc8f76221abc85017edbf8e6d80436a5e61720a508e898697c6c2371d93b814a47c951e2dec4303c93423ce01c98ee41dd2a4fb1c7aaab4b4d7299dadd878b12f5bfc13c678ee0e0fec598724458c4cee8ab604e6828dc8e6d1f85372eed8d4ba402d196f4368944920e7a63def7e41dcfe0092677015d46d86c0264773da4a6d95164463f269523de81cd138fa44eb0c8b34d85eb9c2ecb62b980df64db4c6d6c499e47e932120b560720c0c303a795f358d219c2f362f5842c82a4d0e7dd6616df658586a7bd36fcd4588f7a6e4c727ab29a4c0f556419cb09cf017d1b38a5ea1239deace676ca5006c560972b06e57e58de941c825c297bf2a3bd331359a5390ceff91eecad9b4ed94268b4e7c8720b0bdabddf6a2df752b5e7779e38e12237c5405a945924b4bce6c4a9467c404711fc0c19373d8197ba1906841c9b0896dc6a178eaa81d4d5133b81ddbc2ac9d40230a1a8811990fbcab100b6b72f4d6c94d08d19d448959c65fc6475b59d05cf26e5acd5a557cc0efedea97911be44212482a6d6e1a2987088b49f41e3fcf5c209fc853a5fa2153aaabd682e385e150cd2a78727f8f24f5f2ab1d9bcb2594f4e95c7cf8603bd6f949aed4681af2ad2b6dbbdaa89f1679fe2c537d6594aadc79e8cc290a26bfed7f04ec4ddb84bd40c2372505498ac3d934173f743609de47986694d55948631d0d1bbdd8f6b288d7ca700acd43acf58fc624b570d466cdeae3a122aed1bc37ccd1d567752c1816209087fa33e50fbb9ce25bfa46d9e34eb1386a9637eb0af876693df8540f115b9ebaa9dc012e02733d22d95d998063bafe9dd3a635119757aabbe3cf50961cd7b19d52c59371c42f05b08f45286269f16160c40236958d5868a30e6535bd87311e1afc8539aa8cae1d95b9888ae9f2cdebcb6cfc0feddff96a5219bbc47c5e5dca1e9af4e8119c3c0c4195a842dd5f6bcdca5e37b62632793825647268aafd8ec1fa701a7ed21cf8afba98b9cd098a736224f847f5e93cb4ad107f0f7703fd0b874c85ab21521c252b547e8536c088fee4d0f546c27b1b11cf9a2017ceb49d2b9e0ac7e77c7d57ff196b583de38de2800062a756b9efa9f77a965372c1e839d9d3324d58b4d99c5b89fa9b4ed07103b64b9d49e80f9c9f1da2349c687640f0b87ef32fcd8c6edf32c7c543111b3050fe354b56208519a716dc50d9067a6d6029bfd0f4caaad96a556054fcbd3c5cafff94b994857a12b01ca005581a8627db4cd1df99e1956b49fba3ed806438f7793bb3d54373b00510ca2c2cae760c6dfa93e30725e875cab55af1d49ba3ee5e04fcba7ff9557c50ede5002327bf8e82a1a4d1437f0db183c03a2b52360fbb0a836846cde80f3bbaa656ae915e4cd3fbf4b2bda347ad5b0adbffd13404e1075118e9b6de13563aa895fbcef2f3318c416d0441b671565321be;
    localparam CH_1 = 10000'h45a652e6f1f62085c38a1068a0973c1d214c8ebb67b121a29ca7c6500ff5ec5a851b9f88e88bc2289d420cac4e16871b01d3aad00d86fd14e51f7e26e1239bb261ceb7e16a2b057e758498245d1062b756ff137fe58342911544edfee2674f09f4f1b335c6119ed37b3bcf3af326a513c834609a104e9df40655bd6dc39706c8cdfbc35231292e198b0711045f03a4752f14368c67bf594b49f4d24c90746efccb7b751221b2275ae8c6afda489a147edc06b3b593d5cf09aff8b3e9d90145e70bfadea19f7e8993854d2f542c0f1f25dd5ce4320db494dae5d4851246fa497992fe4105429e997c07357bf6e2a914c207d113fbd84b335b65549a0459a94e2faa941506e6602ba0ec906811476f1aff404d124c79a8e42945af7a65f6ff9fd3001f52089603ed6dc4e440a1df824e0dd63cb90e1427f92b3ecdb65b9bcddc8eb93d2b5a753c06a50ed2fd1617089981af4c6da9a76c22e232bd14a0ba2509f49b68adce7d49fa8ca3aedec474b057b012b9cbf0ea6760f1e7138ed3854504092fd4b483ee3ac98a4c251044d9565f3066f68d81b073883935d3e01d73dfc5f331d585a6ba452f86a01cd9b3cf00cde72408711d001efb953885b02c9dfb0657a10b2b80d9c67cd784212e05ff27467d8f13bc843325cf3f34a59b78d1b99d2d9e132839e5e7ae42840444a5e58a994a617e7bd87d4490db618e865285daa752741aecf45db2ef3a7f953c8afba64e9d97147fc3fc2fd2a010ced24480d3c0318dac14574722aea4696ffb54ea05dbd89f63a8b41440fe30462b0b6a3ce99d2a528f5f046982650e67c0ef929121567467f22b53415ffe4633a87cdfcea914a428db24aa86957d04fec6ae1abd61dced3d402dad536a58630a983ee2c961c7cddc6e1c0d568f804546cf82294a150768b2b013095421ca59cf40b2f650c5bb85cd90c5f6a7097a06d0163fae5a7abb3cd497321fc0742e33b78f848e29fe3b208f932a605d819dcc5d3c09196453512c8228fde8ec85d3d568e5d597e93e572066567d4b717a8e679822027c7f592fcf8c722b6c7e6db2b4bfc9a4e22cee49db6bcf6a72fe8e292f037bafe5e481998b1dfc916b7969b781baef5552c8c6aceaced2c7a188a8136972e7febd451dc85a0edb0d04fc9a2239e05d0813c62066eca3f0ef4ffb36bf17d30ec1ef4eafb60a1cf9f7decd2bbebd8ef00c70950c547e555f02dff66e32a79f372688d4c8b04d9b84e7f4fc3d580482d60a753970e47303dc1e46457548b570fc792834c9d583727e509795eb656f68b37486a2c6b53d74ed183e0506ee7999c2f29771dc6fc5e0da7a72051ec5237e264985225a1da1be5fa0455c257ba308e2b124e6910c1cc2382b4044ec38dda78b74b6829d21be362ea81f2f8fd58f63a1f409d37d99d56306a9fbdcac571eb1cb4b5927f8df121fdc7886ac3adeb43db5f2df50bd4ed41287ff682e0fa93405672983ca4b579d3cfad7a8bdbec5af5857f11a3351ab82aa621a31b9e44b61526fbd27250639c88a1ff0fa86c8092ff2f243beb1bff107d5e4324e27fd5c2be680fbd79094ac4df249242a9beab3df45f4db83117c8ef5c296cce5647f64b17ea4dea3cd21dfd906f18168acf85a93e8fa41ba8b0e790989147e688a0199b0bd4352165295f585560c59698843dba92e48d870a4645c0d9bfb00a5983ceba81a2d5dd3459063a9b5694feccac6671b6cdcd6954fb32069352b7896f589aa8931eb4ed00d8382cb33fa;
    localparam CH_2 = 10000'h442f2f822be27d4b0152c0cbd3c0f8fedea00e23b2088e8cc499ccfa96d8dd99de54d5a58e3c020756ffb05e1d99cc11f75ddff12bff3d9cb6b61d06aa72b904a7d65f8e92ae1c89cc5cb46f502ef2ccf343a548ff5f7cb6b950b2294871aad0e3e36e9cceeadbe23ff97c6c7e0a43939f0d8913191cb28ccc0858bd424ee622908a6b1414071bfe434b82dd73b221d410702f2657a8ffb581fbdc55ad0b411a59aa537fcda1786bfbecbf5da02c1e37a8966c021bb1f78e823ba91736572ef79411c439769cebfbf813d580d52f09a0afd3dbc01ea2b97d2bbf79105339e00d4c7f9890c2aeb7e90bcbbd31dfcee153a49a64b7a3e88a046a2ef774e3de5c8cb6bd8cea307fe142155f8140b779f48ba11b11fe0301add504a93b97ca731d12899a359191d8b44c0a966fd6a57551a151f5cdd34e4c0322984865da72d984743f6c6429016fdbab3ce45101525c043e82727840416ea915b916a4dea9f7709630ac4ed23cefab697b7a5731aaa766be484bd6c32e94e25866a969c52a14588ff3912b55c62ee5d9e0e23b63ee14f05d515142aaddb04e3e27402389d8eddbb0c6ec5d6e477e184d9955268fef233e38b0f474dcee595fd8d281dad0eb96f6317d0b0fb62cdd3708667d1a4b42da8b6263e12196502f7adba6d46c665b6351644c4eff54bea76c68d13492c858d633423ead22886b525e6e75805ad7ec3222e49f76cf953a18205b16535dba26c8d62abdbcb64d295ef982ee080af1a86ab8389298035e9a5528aafadb040b8b72df951447c79226804be05367f65c9942fc532172c4b6b3e9f06dd768171e84c3d2c890a83cc3b935535d48729922e5b931f432f0d94ae2e8af18e5cd172a8a2c2fa4d04bb1645c764e70ca901e814d3ac1be7403f89600b059adce7a5683c4dcac041b7a57ddb52678ad9577383404ece94f7fa195f36cd99f0889e93b00cd75eaced2f08733ad4006adbbeacc7a26c5e66e1f33afd42470f5257c1f289d6656e813ad0f9a8d18f5b6ce6ea44c814c46e20d57695f4a9436eaf2a5afa6a1f72c62df98257f79588213226e978f095f49f02e682726748c98edb4d0661ebf52852d77a2538eb0d2615ea63bc727e1aaa0df0e41dcf0826c977fd116b4a466f676a02372c75abb506c1efb8845857f9a4a6b1dc21c11f45431c07aa69d8fdad0348e0e785c8b5acee8517ce589d3723e785a6b80d00cd15dd880976c15ca1b58a8dff30262bdd84d9b4c0c688b0b4d510565b83235bfa78574a5c50ade58b552fae0ff616b486b53e6c2d44b34e3b2ce3ea977db870c9f8759dd22cd99950752cf2b8c229be82325b75fc4dec129afcc0960656cfd561f1142ef2e16c76b807505eaf4de4fadc0d268efa642e0f86f3dafc939617d103e2d99419703b48d4a74b96a5886e40474beca5874664f2492865c39550ff8c1133c81636cd9cecef5c92490e1b12756c0581bcf4e1a71be4dd30d64b743d2645d842d6c6b8b6448eb51162c776c47d59f471a20a3fa69a7361458f20087ebdc94de676e717687642fe7f59933164cec0aa787d33e5fda595e2e325ab733bd04dda238a6bc050e31372064054be58f1a323a1179839be0eb1cbbfe750cd5916f3c9e8ec80109dc9ece57aeecee21660404a8e3e334fd212d950ad548442b0b412888df9820b552066c2aacfb8af2db50ac2a5e4159d1b7c92e318b33de233179fe682e8511ad6a30550b5c3caae9eef5566519d302b7fe578fc77fd74794e5;
    localparam CH_3 = 10000'h93a5e7159b48e7c00b8c058f5d0a5126698db08eac4bcdf54592ca294cf8f9d2971deec7cbba924975526e735151bbc38ec00aff6c8dedebb80d7fe28aba5aea606c591474738624156b5e73389873d2a6c7165d5b9b1a4c0f01053d91217a419be5e8d44f2125a126be65d3452bc37f0b486dee87e3c11503951f403cf4b20324248fe215f85abcec27307c9a4c1b71a8a8c5242d3612a1e85fec57e9e003601e74e924166e75e66b87b930377f348480e1a9499e37aa9af603aa325e59a5f8ede54d1273f221a0185eb96dff176094370ebdf42c21caef57ba687d45003fc0e253283a956bbc3cb059b149d4f8cd670e6992ceef3575330e6aa798910dc4e21c38ef0800f5eab4f8c2d337f0022dea6e26df4ae386b4eb0f17cfedaae990e4524a8eb7dfe42affa48eae566118977a7d7ce42cc68ba126d49b97cee4ffcc6d0a5927fec68a534b1294e02b97e2f68f9eee3c365aac4b648b3711f8e272612df1b286ccde60321c070cf0ff2aa493ed6b916690dc16ba5392eb666d32bf653e1aab26809c992a082439ae69e0f1fb4dd9eb4e05d3f475fa6641ffa65a3843cdece485a386dfba9982c38f562f21d73e1df00e9b0ad5099bed7dbe1c185139dc1f23e9fb7a2f51f22d1ab68081d92415a460df36b87647cc85cfd37bd5972155025a68d82a032b66cddb8315b3f7526303c5897a45be1f2cfeb096d50b72333f52c21f6a6826275f365fb09e9bd6f2ed567a97b6e243b68381c9446c337587f436544d93c4d83e7c5f2b4d9460ad799372d3cb957a80f436e53fc179e9ca6ed1280b34cfde484bcc62bd13e4319d4248cba61107920ffe12383391c899747c2f4e176b409d409739720e842229b5068b0a797261b9a3fd3df27cef36c3c600675db69bbf9ec6f2730b1951d88f20501deccb873ca0d7c4873d3e5f991cb3154fe0b2834ee0b1a4773f64e9205706fe554997aefd9a9d7d475adf9674970f60d7b4f4810e04f5e64e529e8736f3b6527298048510274dd9eee740ba3859ebf6de0e616bff6664efbc060b61959d76248f7dd8f5c5f7db713fe17efaa094afc24bc2aa65e9aa148c1a5207701ab2df7fecfac337548b9b1eea930e31d76bd9bd3d31fc82ba9bcc5faedcf19b72eddb61af20a7367205f5e034d538f1d1b94c89fdca5498a526252d1599f0dc66d286424c086a1403cb225ea46ca608630c6cf5a1841f5efaf2e024b84847a00d24bd3e58535aef49354c0dd011841fa035dc973fcb5f6d600acfc5055b5b5c9bdb7e60dfa2fb887689c90cc22954ab8582429d51772a44ee68a1f254782fe65c12973b0b956da92cf716ca17ff71d5306b9b27f5664354ef52059ae4544e651273a349914875f0fc4600d1548efb069e8dbbee8a5e95a564ee81aef6b2da9de64712c4a40306fd169129d70b4ef51403b2620a15fd917d79ba92a686b4744d8d45ede078876a975bc395a4382b25c3f5445ab8b30c23422382f29f951d0729f1917607b8b4ba1d82c628712c8876baf0c48c811bd42a700e85524712dc47badbfef6812acd734ea5de72f4b7106e22c23076579ad03ea13061a4cb7ffbc9bfb0c97d8c9894f82e6dd5ea32d642d653300eb85d9e010b228d2f216cb5131e6abde6fa52beb2a9fbc0157b24d57cca7353d954c39aa3a7b69132509675f9df51a272acf4574d58f022084c2a4907143223c4129b55a2a28f7f8250822e2409127690483ec265c18332e0653bd99a58827cbc8b8544cb8;
    localparam CH_4 = 10000'hbcde0061e457d522a8f2e2ed66c59875629f249992ba17e1f23de55dc0c9dbee1d56f650506adf762cd09957f1a19607732987312c648390b38337be41f6c6cd79df8d20efcc044db7c625118e3a3c835517288b1053b6fa1d777b4d2b0e06ddd5d96f36c7bc63bb89b30ccad0ed89531ca9e649612a2189473b29dad43955ba8159ba016163b10e7a7e911f120553556fc534816686d61c01408a3492979c99b5d4adba2ce8fbbacc1dcb17cc948f405dfa8d1e23c6585cb0376be5fdaa13d18183037c14b157bbbc29908d9e976e1cc4ef62ba50431537b7a593c0a5d890ca240290ae1809694b8797904bc334944aa4de90423e6416e9a592bffd476781e7a8d21f96c539cee1c275ff0fb054097a1c07882535fe7c19b799cd51f96c346fad1305c19e6894f89ebe081f898dc7f7adc0942a48d9856478686c04f70ff6f8cdbfda09fa5b6225a5ca7c2aab42579647064ea8cb097d1dd7c40136b61a85dce130bb402f83eceb7e90b15210446a8fa0dd620f7dd59bb868f1c37ec5026f89087acac8ff07f74b1d4d043cd45e9ff3f5776cc10e88e8eb4f2d34bc7a50ef6c4caf571a8a96c656447b72a511f950b6e84f4506088e32105cbf98b59bd6b0bda0dda2eb5bda5d0972482589233dc1d5b13ccf235c7b3b48601382487badef8a3cd81a377d58d49f35481bf9544a04a284c61a5a110610b5b8a185494f547661c4536d244bcf2d528f0a1a71538cb218e047e0cbbe5a6f7ef31b2ebbc5af906e087a039f460b3a9bdd5ddfce96991e0f31121be83771107f7995009a9b63eac04840cdf48bc060c756dd8b41be94c40a1b8fc935765c5aac479a9f9b08c9440260da98b088ba031f59bbf138df32480366b1ff6a76e1690d180e268fcde0305774082f18319c50cdbfa0c25a17522c258b99bdfc0aa788515b30def9b1835ff9bd34017b406c42ee28cca9c2b2e5063b65043dd8ef38901fc201b948535837e872e047b19ec75ed8baca32448cea3be576b072f03befff3c8fc98f1e7f04cc174bab2187fb8bfd284115277253bdaa262f1b523f4610d963de62c68c86c9d57ba78b60b8abf6793f4cde7fbd2912da53918c573ff643ff187883062c322f1cd8b4b575fb0d3df6f61a0743579ffd8ef46f60b5525c28d032802a19c9c7b56131c1050931c3f2a9942eea1180fbd0e2f6897da478fa0964815254ce589cef841081b56288c33a09ed6d2e42145a4ef7be3281ac952a206687ced4a2bbba52bc7150ff5196ccf5530363cf2c5b86c62a930b391cf8ccfd9344038157cd106d2524397515755ac5940f8128933f05caae043fde4597904a4ae9eedc61e794c827adf8afef861fd7b16e90869992c984eac1fcdfd56ba7e243b8a7aedc0cbef981d782089778878e91cd563939b0f8a3e4afbb2038b17cde4b54ca70aec942511aa0355ec1bb1a73f94433bf943746b1614cdb591aead61f46a40c3f4667fbbe770b1cde0cf457f91bb98ed47f002f2d4929ac0a89dbe08de3d4be704a1d679e0d98b005f252cedae6b3a546d0006268c4ca1ed8591cd8a898ae13fd153cf7be696e9bf74c39336fb3082adf5ee0816ec7d858c647139270b0feef1ebedd3b4fce88e476f44ef29d98f05917afb5c801f8f75ac50bd200f0c7cbf5a34d860f197966a2a1c6d7ff29b8757672ea2a23e5bf7b52faf2713a098db27a8d7dc5bbe63b38373a286837d3b7ff66fc5001dcfe7bf647b7b6821578c8e8f47cba973bf49742d017;
    localparam CH_5 = 10000'hf50038760b60d1202db22781e2ff66f297c84d77fbe6c9c8a697e7ed468018a21efd1b18fa52cd6fe13208ce8796414a0b9fec3568c86a7ee43e37f7de778cd7f9bdb63a4a70300661afd26a2ce4aba8259cf7565f50172cc52d7c0e677468f790900ef439d00359696258d504ef7ab89361f2bdb02060dac6c96c672db15c2e970cc7e581643cbfbec5c4f9cb6d3ddd165d8c4592243a1f16af07b1bc9c202dac713337828dd3afec76425385a2426e33fe5df5efd66e06faaa615007c0ef3737c087253e979b6c33450b3af8d697624b396a4d9a41dfc65ba838b2092c9e31fd43b2a2beb0ac6d0c39b435b417cc2a0ff432eb06d13c3fb5fb9b5df4fd1f26c30c1f68da054e116c5de807fc7fd56c920e6cb9b20397f73ba5318c756d717740183181067a3fba75596fffe9a9371d545b79f84f1e706e785b8479888cb970eec3fc8b6148d725e4613b5bee63d9042a1a81dbd3f4634b77c9d740a2987751e124d87b7aea6d554011d47a0af47758280560e2fe25c3a6ba699eea102cfae8881097ff76e98954eb55738be55f2d20b219529b1da4768b2025a5981947224e18680df52674c076ce7d6f6eeedf4c33e49f4df7961bde8d8fbbf035158c84e4f4cd3c840b956f28cf63d68c602f8ba928fd8429dc5e88f5824fe46e45add383febafb4629f7358fdb9c3d505ccd52c0ab30703e523fcb35330afc787f5659804767fa1147f6efab365b232441bb44e24dc8f1716fd47c1432e03dc87a568fc279e154109c6de152543110f6f7b67faac9e025714a997be9c6a60866363115c9c4ab01b15d626cce415713b6e5514afd5c760be5f02634df96e8cdb8d5768acd909c95a824fa971833c75451b1cc69651ad00ba6ed4f43ed12b8faf4ede1ababe57717cf524d6888b71ce4ce5566df2689bad812b0c0c061f538630bac1a752c7c19c2377c6c833ebc00827f0fd1ddb5e4708a678fe6a3b849d3f1572d20907a3f023da40c55284b095fd8b5e022fcfc14e042f67f133456482cf0d0961d1b2a5d24e6e823b313a16183b5de4eff2877ed4dbf7fc8932f4f9343089ef90269e3b20dbfac8cf54f6a89f97234d4dca2b14cf8ea19c1464e5feb181e0f4edf335c2e93e91a8383b4bc20c18f232009cac541011a2acfe34d3cfdddeda77c219e8c8a33ae50fc501f7544a79c1250d6f21d242278d3191eb026bd211da6a95f55426531741986f784382f35b1b362fdd5878bcc1583fee1a39843dd2e9833251470b1c151a5b8a8c597fd998e622dec1f4f61e8e6d60a5ea7f9ad40ba1596ad4616339f21d6b136b80a2f81ddb3f5b8f925f08dce9ba184c96236c6b7882ad3baaaf5d8d3dd2db2e32484049611f65081fec3769c0490bc5fd80fe7edb48de03ad29260b06601600775132574cc2008a49bbbc0298f914a3ef6dd36891a54ed60091cdfe29718afba7ee3c83efb571af3f1ddf9eb967e2349830be328f1cec4622347e9502177462b79e49b7b524c8b46bb2308ec3fa9c0f3edae476fd6ea8c16b5b620f43a9bf6aaea1c00c44a536f3e51a93c1f1d19d15630625943767429d8489db1ab855fbb12d701ac4b589f8c7dd15d18d004b9e9e48945efe2200c195bcdc8128ee19392b13398492dd9b36afa03c3bc7d210426715c5adb9535a015518608b85dff4078fbb536700a1527bf0c87a41c8f6c6f1e2b016630cc490063e64be2cdd301d17635a2078174bc52304a2494dc009ce76253b44375635234879046d1cf;
    localparam CH_6 = 10000'ha5f586be4a6a29f0e6377700a5b10f090b1f169d0044a5210290ec61f974dd010062864385aa2e77b28c5c20e83c84271d3a8ad2de9fe75905141db639bcd653e154d1e1bd2a79485e74ec1f18fed205528be009a4c1fa810edf640cb8fb51b547543c8f306975347be4e0ff06607d856dc0ed40073701379aaeadd4887db7084746d7c60ff50ef5927a28dc95d308c0a3c7b4cf99803c5cebfa930c63aac9475defceffdaaec305affef378a49d11727e0a2a9609f1bb92e056f297681918f4277af43533da73f484f8cb44a03f19fd1f398ce1e933400ee771e7ca9197c5cd5ca9ea192c3a2ea51fe135402929b8025931c101e170dd3ab84217e67be0bafe97de3df9b38622e2d43dbfda51fe77e81e12a132a8a0278bbe350e633423823e28bacf0b205749aed4d58251ce0bb1641f162a37633ef9f686bd567f81763b68d7c13098458dc0892a2c02bdde02ab1b4e16b97b66102dff3a83e241ad544ca7860e62f54a7eda7a7ba891dc4becd5c6030a7407d944af1864207731ea12a2580d362b6e5080824dc314c1d0f9d7b587cc19d867a5d7b43476ab78eaee6b6048436c51042d728ad63abfe130dbd79ecdea513fa8ffc243b6374e442d796b80b311526e06ac41ff896640d61912aab9cd556557441497129fba6de991f9d76af1b4b307a6cf67ecf8219ea8b9db87d889abe63dbea6509cdcbbcc872bfcfc0c1109ac3797762d37d5c8dd8e86545c3a651bdb2b083e71ff98d19fc80b5f539c86bd0c0c4ac16e59434c14b04b21aeafc7021033deddd7d7486cb8e3940ae59e4ffcd24dce3fcfe40c960d7f4340c0e5fdfc9c3168515161de9891a18abb81a5b19b555d2b50223437fe964d4f4c42861dd0ab1f576513b2278f32f1af5c76cc40bd91800fff266e0f4d877068f4917cdabd27446703b8f7885786eaedfa18d052bb0c92bf675502cdb4935ef453ee8ee1a3a8a2358c665ed898f8b8af0c751e76753fe31dd2ee464b8baf747a1a6e039cfe6d9c1fd14a00bb01a4b34aecd90b7932e7f206cf51aea631043f8b54aa83f6b90aeefc85e026dc3ad92382d12ee290dd992d542cc0408d6af980ed10c9b5555e954fc7fda29236dd54e96a8be23ea1f4816b885b8f4b019d7302e5a3b895b7a11b92af38e5ca50ed301a12b295ee2998aff656ed25084b132704bbaa71ca9cb1172d59b19de4a222c93fd833bf907bc088bf876bfa66b7f129b88e9e442cd3431f7692d1381cb129867584fc36fb4d3e26d8d6f4e6d52078ca04d6cb96ae81e413a86478394cfea177be0fa6031307ca7d89204bddc3dc18402b59fa2ad179f0222f3bc361744911efe91ed5bbeca8c0e4185c1243eb5e5f302b17a7243f726489d3a747319cedb534234fb3161fa13055fb00a4772e9b370a9a0917e5538a5d950f2d01c6e543b41797853448fa1f9dac74f7f6d3a4d9067efa6e9e4612d8a759cc01161de1b5ddf4b0739fabe27a715944fc16592a7c5b6d5eb15ad616505e28c6b4e6b94c89278f8d45446fc47ec40809c0da9ea5fee745cc5b57b6f282c14d5d2953792a43a99929cdca75b53722356db0b49562a9a52cd3806b8b98746ed0afd893e5a95b734e1b195545c614b6db78de8586f0282f09de607c723e32aa980bcc542c5f01e678cf7957bd0cd4c576609795b20e4f4f4095b9bde215523c7be2ae5dce34433e45896a88464a165c584fbca6350cafda1b8b45c58fe75ba446056dd5ef5e49af2a43d2b162db4c3863;
    localparam CH_7 = 10000'h14045fba66beb079cda03d4dd9571afa48eb2904dba52c121f5bee66907aa7d7938393de0d7ad453711e881fb73a65520b1e130db95a99dab4a017f9d9df971d4c492b73d08d80e7e476402ea71942d55b6f35676de3103fe7613d3ec350e740668640e6d8d39bc6c2cbf45319ee859f80559cb1ebe504b7e2c289b4360369a0febc6f148d54a067c56d55546ffdd3a7ef0ea13ee0a47e341e37dc05ae041ddf0a04638de9232f20757ecaf8edbae10c910cdc6e4f424ad35cc8c180bd1a0afe0b21ed0887dbba233b5d75a867fb73fe43f1bda841a20ddd9173648194a53073e425e62e60eb601e946c8aa0e975995d5504d1e706a613fbd744da6169212954b7268d1817a12d0d21e70c3e9bf334cc0c7f954f6d7732d6bd0f480404a515dcc69973bddcb933c9a8e29b6e28205cfca64eaf27ccc1a877c94b333767f69321c39b80071f9d579078f1a90d56d41d4bdcc07a8a690733e1d00600601495a74fb1250e68b6795b3a7cc984c591996ff688a3bd430050f14e1c337aa73d0302c745eac9207f272ff2f3ee943e2721bcedd9e7938d6019aefafb9e9630876bb1fcf14b9a3ecc577e02dd325e81ecf0b618fb41b20ee8cb9ef6eafd3637de0280881e91897adea4f81e9469b9b3552c224aa4c13ef8aeb9de1d6ff12448e6dcb38b124a1c45ff688d1e27530b13eb7af96bafa294d00b97c18cecaa47974cb3716b972193bd57fa2acf83865a88939394437d1fe560a2de60c78c8a59e1e33695d199eed361eaab079b18538432496f42f490f53eb8c12d59e2aee45eea3abf18b11cd333e092a01a93bfdca84c03bbf7301dfc8dd640b1f7999faaf5156f7c4417ad55b331d2c99508d35156f23472ae83ec08eaa57dc52f7acc2f21aac5c6cba2923128ece7798b45aed46277a9883a24f032e3e415477059efd4ab3d9ddb5ddd7047230e7b9e57b14c302018f181d0d7c622c1af92097a2355196dd915ccba10baee5f93fbf240905c26b04fc157f5228d41e4da4081408e77fd194dde673d567e9e494c0e58cacc8a1e339b53003021a1662bb4e174c50adb4daa20e5688512841b7a67f92b835e904e2e74ac41b6a74776ee2ea75029b8ced9c7149ede7dd0e848e2e45e0fb4215418c26b443abb05cad7ec27e1bf41d0a34920179aed529bafb1e888f0d18c885ddb210abba887fa9e3a7b64b6af3f948694de4d076e606069783b670e5198494e8699a02848370d6280c54a80b6e24ac0cb5ad286ed673e030dfdb6b1ecab5e0e1c78ed9566ae4e4c79451f52f372b34afdc76fda7b8c97562a31327ec8a3baaa9f12fb1a6f6502e10246aca71d18b6c05a83a0570cc2d31f08ad99ea989de2b963b05e3cb78efc2179b66152219826cd6a57e54b11bf74890b27de91b4bf746700cd0b80c2c35a77a95fe0d1209b62442841e738e568c9663343d8eded8078a636e59a0bfb5dc2746620137ed19a1ee0710849a2c6ce8bee77fb4eab4eb10203a63f35aea150035ad32a19cb97b3521f3e8671a774fb529ec0aa9cecbafef2d01f57f1f52b8453cce857f2bb29d2520de5922be99a0c62113a827edba0afefae48db924f1ed385e97573fd29568ab2a8ebf3fefdf1a6690840df34a220609536d180af04cec8c1f6d4a87a78fdf85064a441072fe9fa26e49d1cabf47ac2394bb838af75e356bd4860ec4311c085ebd7c7f6e00bdef79d4f7b4b7608ca8865d85f10b8b06dd1d6899aff74501e496de7b545ee2a0392e45500;
    localparam CH_8 = 10000'h8146ebd508faa9c38569c7bbaba43868bef81c38e4133ed6cef4c94cfe2d99ec1bfdd0bae0ece1495d6718eade57160f31e926c4f6065ba1fee48a611d35bd1d96f989a6b297184915cb8d14318e9782770a327e5f27966e99b1742641806d909209df58e66590fcbc391587e4ef72dbc19e1f6f13501cce4baa6c00ab928d8890af59f0c033c0032805796315ea4d52113d19b7b8c095aa968d298254fb58151fe9f7f7e036e776374213442731b525207a7d725346b6c531db1d75e523ea149c16102380d4e71d1675f94188c552baea10a754d4520440a4506f366bce31026601506b23981a19cb9bf14cf3dddf69e1103b3b5c791f2a57d882ae3bd7f09b8dd1002a8b2f743406cc6c2fd7d2d7ec39cf017e0fe89eadc2caf184dc118475d422c35ef3985d2f8aa536f8f97699673f9ff3f806f5c3a463452fa000f7a21aa592a7555f549c4e6d2ddf63e9f21d7bdd98c2da9dfedd0c0bb0f11fa50173b7135bb3e6143a127a03a76b0570ee3b255eb17937c20826e2e54efc13c9b1b8a24b4c5113da15a3edace96d64f2ecd1fe77e8750a92f6817c4d8870ab5d8fb592020e385e69d31c7fc2584e05b7bbd88ce59c1a8d1a4e17ddf247919fedf0d4e0229d5de445b2f30a5ade4cfabba7f10a0c01ef9a9cdd8207e7ef3eec7361a6c07dc25aad9f4db8b3646f1aa9ef23583ec64af42856813ee0e8bc6594f490d5a82d055b6dc3032d4d2136ce8611f52f9bd462ee04a24b79f0fe4ad38993e06842152ee9dd48700358604674bb06a420e42eefd41c5d4d35f9290485a3a84cb9fffb95412f916c57caf845d337c83d7f617dab616deea6aa6d374e1cdf768b34b1eb5ebf01210377d0111ba594fbcdc21e713e362a73228b5617f1257a5ba4113d29b609569e0e157806721a01f812cff4bdb3959e308812b622f9d1db7af2a2b97b564c5bbdf470963cd2ae20538500fe933ee7e3bfd251a6769c04fec717517c69d9f4cde621f97632437bfe9bf4458b3368b72bd3b383769f3c881cf007e6ddc9b48d14e4ec242b12e2c127b658a89dc9889365eaa8dbf8714738a4150c5e7edbcb52b3673f6ef16c0f9c8b35ca8499992101d34c0a943ac50da7b55fe026b26669bff945f9fcf64800d6fc420d0a506726fc62386604c21f13f903184cb450e6a30740fb5150757e37c1eb4553da2d9200bbe370ae78cb6b754adf591d9d0d2ec49490e0468e331fe89f62cfed64e42cfa67a2197a4f07e7bffdf04c010e59823e33c1cd42c96c368559074e7cb36995f2fe920ee317bd7d2fbd84f9f38d41bd1b02f26a8a20c46e61ac51ef22c5bd1628dcf5c7caca55808d655d8326777016cc6c25c0f803658b3a498e32d8ca02e9e9a9ae9144e13b81f09f2c3adde33f5ab2425835f3f95467fabcf51c187962390e4b9484a065df0a4f40ab0ee58d0b17aacb190749a773535cb83ac44ec21f56c4e0d3e3fb80207252a06a954efa3bd0041d23fce8a3d7c969184a39fa8a1aa367d1f0fa28efeea18d8787cc4e02ad77269954ad3d43befa67925d1c25ffb714aa1152bb1e305165a2b89de9fe9b021d2a97b3fb0574f22f26087fb8d9c435b183d3c095b666a10b001a3681a94aac0499c0b41c57e05b1f4b40991c3b62a426e0cd59d41506cf98f5056edcf8ba7c19d522bc1e7beefe1877bc17aaf8394c9a3d4420d03a4ab253bf1f2e55b35fab9a617d04a69fa000b03eba6e20af3dda92e46037a3e03f2fc868a006125aaabb69d7;
    localparam CH_9 = 10000'hfb51967a1c0efa08326bcd60cf2bdecc2848a8b950f8e8af95220175201eaed7f485f0eb21f89250e4bb317f08771d17c9749d79e009cc94456fa2c4c1c29f504daf999f492faca34d0309f2780411361dcbb80f0c32e96bca394dbae7d8e4c22cb3a49b880e0a9dc2af322f8c1bef4e30538e7c6752a4afbe69e7116fcfeebaa0ce1c700453cf028a86ee96dbeb8f82f6fb50b870da9437c62013f1a78ce4c2bf0a85958f0af75194a8d57b04aac894e71d542ba71104963d2235289ad20e0dab07f8af949716f713c4bd97f298ed12a2735ca5503719b3b9b0b6fb6a34498207cdba36d05fcdc69371371ecfc41c1a073a427734373f758f564b85337bd3d80cfcf01961c3a56b61187379068c5bb4035079ce88196c34564c3185d9fb93e21f4c707a738650fa80d3aa3ab1b9924e341276d3cb3335bfd80cd30616df4e5cca7c80dca9b3b1276e96ac19d724ea4c8dc4cb36e5172fc7de60d3b7235982bcc83eee1158961b90cf033da43afc844791ba274f2c8442792b04dc139016c44a1fde23b2d8cdc2f5eea64c276d34591785d00448a4a95bb48dd90e0d35a07344f21eaf42239e07347e77c6e89c37e921ea6caa8776a3bff903c14a90f48244c8e4b00ce017bf04266a858dc805541ada8f6ab5ecd46acae5e63a5179e0e29329ea9276bc8e8d6ceb910f09a021dca40cc571b1916d8f56ad57bb9d6f0b0c220e1e79b0a7f9e0bdd1f2f75ff5ae054a786a7b77ce983a192e2f762e782909358a185c253539f8ff4394843ce7fbf6bb9224e03fbea351a104dd95e1149bb8b51b7121c753b0f688aee4b131aae958011e9d45e33b95ab57e30801b5e82c2cabd6afd1a39e9d0f3a1fcfb9d10bfae1e4918354affba6630a05d9f80f562d2bd1b3fa3a851e416ac8e3ecdc1fdf7e9a099b304e46e6ed1e3d4fe545a17f62c742b2c1531644ac701d73c47ff53adf9a62b4aa4abeb9440f4c1270562c9d37f950d66c69a90084fd38f21d7ffc25c4059c2f52b761c554130eff516aa24e7edf67fa5263bb52dfd9a93d1caede80714b2be5117ecb03124f8a219cef998435af3f18bcdb11d885690a07814f254cc03d7f4176d98a93fdfd99b65eca79ef92e8fb36b8f656fdabe9c514c07170c41ac6da418011c550bd6f0f7ed9f053f1e35b43fa728723eab71b48b3cb5b70c29867e6354ec63a7aaf73a7aae5df7c0902210af54112d990f51ed58ba6ea201c3d469ed67b76f0ecd97c085093ed69a8aebc16733c3315609763c211d2be4339eb807be08db8cc983bcf288e7cfe792cb3cd00d68ac2df08613f746c5d6c3220d1caad786debb8b7a661d83b7dc93c59f62773631dbe583563c1f29928c698052bb8e7e509558d408e5929e2b7dcd2b88c08981a31ccfa6ce6f4e0e1c3d793abc61be5283fca398015ca1b00f58ac3a752cd1e924022954a4b2e5853f03d5fc58f8c2604be2a9ee3a3c18f9343906fbb14215b9ddb0d98b77d934dc7f6a87ae7905165835b637f3397d50dd9487befb8cff42f3f64019299c42e86588e1092f11148358fac39330c2c951fb9bad26f720b7515df58c167a4ebb369d04f13a9302e8133b664f6755d3aebc56f2425f3643c69f01015b20d582d2f4524784697054bfcdc17911e637bc7fe25ca5ac584889178dc870a107a8aea9ad17bf53136ec32463cc73780245086aa42737ae7b825df6dae608a5171e1cf77bfe84e86ea03cdbc82a34cb46aec300811dc830dca0c0df25d75d741;
    localparam CH_10 = 10000'he229b78f9d0f3832023caf523b1406c78698611a0a62cfafb777e14ee5e27c67983d88fbef42346345519826cbf257fa7479f865a85c5a0a98924c9d39bb6befa83a421b32a4fd6204633f7f407d9bc0abe8e0d65cf499ff80bc526bc3d6427b48ca0e6e231dd335f7eb4c544b8920a177a0a24f8ad0e2c4c9fd6ca401e65f53d2acbb347c01939bd2f62c0b85aaefc86a35e5dabc2f7dbb03c2438ad51ff65bfb66dd4071a1479cd0d88a658ac246f03486bef570a8718b6622d840243a0904e8c2504be0525f44ffa17608a0660faa591308f80c3c6e47eff028100c4b071cfc0d9fed1a1470c32fb0d1e8f0bc47b51aa9e933a9b31864efe81d471cc486b4da0c4b1b23667ae81cafa6f66f239829937beac69e1b9d6e1568bb3c7ce11125b2e1ecebfb6cc63b4ae375c8fb7d5c3844581dbe0765be29008545dd614f893591d45ee4d7964ee081744d300fb29961b14038be330750ec4f47ec4ad5ef34868969560e52c64a154fa0518565bdeae0db7aefa252d56017815a3540508ee3f95d2f49751a64595d292c675fe13cba4d709ca229e3736ac8a9041c5baddbab21ddedb035c90f95d0d5852b025ca4d289cf6792dfe90ec7987397bcadb6ea2de6adf8fb7d7b33d6add768879bbbb2cd2ff71b0acb17fdf36915c60475f9812d17aceb4c4534e3f3590990cc07bff0793a691f846ece22b350881220f75b1d7c6c1258c3a4b7370a9f91b61c0782b39f23c89219edfaa2531efbda9d597d9fbd7eace5f4291b2ae8eb191d82e791e355444c0f8e8826298e57569ac6438c6dcb534b5cdd72cd6a07f192568c7e39e0fcfbd3fdf1a98db0051b14d0050ac9b60e4acaa9ba75eca44f6c9a48fd6d77f00d454de1ab62c31b977e238bd90f79f59730a4e62590d38097fb6359741c00baaf8e4465115b4cf3fe3220985f38b93063c3bb5fb1b2a520b7f18f94c3819bdbaacead5ea6bb8b5aff7b786a874d294337f7cf750af40bef4f39ce606db964722ea6edb974892f3ac3d4e8ea0287fd992acaf0a4f40dc2b5d844abf393f6d3c25b44a93f414e2d4158fc46d2da241bbded4eaa049ef976cc9cdbae27067c54f076262fad1ad93158a2a4502f665a87f918ec9c1346f36dde451dc074369dc5ba97630eb875aae0b66abffcb715ecad59712313ae879c124c77d56c863281956a20fe21ac0b0b22a9bd944c6bab85ab2f2ec8ad02a98d29cb2fd5ea9a1bf57e804ede1c1f504c86e0dc82f3fa70babf4b485ff8c492c8aeef3386cd5bb75188c423477bf17c29197af65497e0c76c163dbbff5f32d568e51a3edbcf374dba2062e85bd6c2015b36f07f418c8708e7381a20977b54dd7c5ff052e694e480839f7ff136588a9905e3341121b476a85f66bc52c370a6f9d553ed8dc9bef20d7302f4e804a874dd94d78c456c111f550e78f49e86c618995156f290389d7ba80dea2681f832808132423002db9b5e0fbf8122709565b1e9d263572dbc5287f4030669195c4ab1111ebd4391df6869b1d4ce45a92fb503df4c906d2688310e9899f9bdf200004aa9a1f3224b414808fbe151566782b61a8a9b23a183c9d9168fa01e550d21efa1abb60da25b6a44e7d1183b932663f1747329fe02269c1284840e64bb5a097e75b85d90f5e0c0d21090e647dfe57d7e06bdbe38a9df03a9f54fd51f58932e43f6c262ae6a7e286c3c7120785a6652abb207f9bd14c91218adc905b1f981902014d00c03ac01b107a82cdd6fa1d23a738a;
    localparam CH_11 = 10000'h4c0334fdc20154ed1958041f37ded872853f73f322a9a1f416f3bfbd0e92582fb0388c44506465440d4baf386a91faf5fe7a70d259261173e38eaf1f3509e820ca1ff087312d4ded08550d3c20289093bc9a3c6bba3fba6817474785fee09dcc46e3566f849fbe475af34cf805efd33fcabc1091f3ed69b1885ef935a554cd012d4de3f3795a625835e857fdff6dc1a0f4840cdd6aed369ec490b78ddc0dbd57fa1d6ed7c03391c5d6b9e17ebfc1e5979ff7a235a082e4a67623aaa22cf01f1c34710370ccece0a82cbde6a39c226b15dc9d6d53d9365b830496965ff613919b645385cd76665b7868fac751505468c7bb7d08284284cc9033c63d853e3f5e14a7c141971d93ef8bf5d240ed12b2426a4b5d3783f87fef832fcb04779ee6a5ba9c12dab86e39216552d2922d9144aa4f47271baba1ba1b9058f4e92674a1102761741b60c2d1e389e4d005ab085613cae54c452574f92ae15ae12051b8d9e4fabb1e385655d1670d7b86a14105e481a4daef5fc0f0609cf486e8f5b18cdc6f117add54e937782baae4279fcf14dbe7d22d09aac39113c413d6511ac47a6965faeae86846fdc0c1a49fd8f884335b3e2ee5525b377b05fac0185b9a2d539a7ebe537b0e793a33f0b68b802897f2f5d32e0a11f9f7a5481ceb91cf0aefc412d7726a6d4f25ac144718c31ef6c58a12b3631b7cfc3d8fdfab59b63e14bf6f17529643c7844b00e7e1affd229c8ac9de7bcf78ba1b6c9881a136a56e7ffffefc9f8424e903c5eba010beb790b1a06137a45c645dda88f9b52151b16c422a440bcbe52e7d9b23905d0304cee2a571596dbf2de82d7c0b50603647a3cf025fd21d63c16305b2fa3019f9632902306fdb4c629ab1d2ffd53eba80ee9489d36bc673c7b74babe29921db403d531efcff37c66e7d5d4b3a580fd0fa26bfe3e18c51b4105a1737935a6919e2c3de15131cce31d23eb1556470c994bbf7e5b4f9ccf55b484700fa80dd1c5ecd77556c68e48cfbd20c591d7fdf556ca83008407e6a22b310c4516d9e7b271cf851b621fac0cd2a010c3e3e6034983adfc1ae0aa58e19af55c7129a890b0cdcf948bfcaafd81759ba75ecdf5a6218c27f4dae604f7d20a3c6b7f43f761672b05dc3b38285b21149574c4c03a947ba9f7a7105036cccb2ac231dd9ec0f0c1e122c0c3ca04ec0de9ee8bfb8f2daf090688341d841a42dba1d65dae13de8644e35dae82337926299fb9896029943658d3d9814962c5d720fef55006ea73e9e45d61f84acce5a0f0f49f7147e058a4735dee80eeae61a78e0e349d65dc463e94589c2d2db2bc76145b5472d2781da2e91c6e4c8c87e14344f062b01d16eec0f7b693011cc4d7b4c3457cf334b349abe9f9e7b4afe840f6cae2129cc89f082bfbeb6972a26afd33701b38c7832de74df091e07c5a773ba7a562c811acabfbc6ee4187ac8d32a41a9f4c12f4d1b2647508d2318894435dc65282c23adf1eec7c40290af8a2d6e69083bd8a52dad7862b6b30a0f0f4863f26aaaf1d7ade94d0e8e9f00db026db764949c56f6f5930c58dbda3ba7059a0948eff842fe19b4fa1c4630a7c83a2b22b4d39721827a747c3e6b27045e5f03769109998318678ef097d18fcac0405080fe331bdb594dbb484208f5cf0bdb2f94a563ce0c4b7a7121ca67e4379340e87245fcf7a5492071318bba41f300f59ce0de37542af39548ea7ae9eedd8d1d69e5d8f5346e16168ac3f2219d8c50fb825a2122b3b2a4153910;
    localparam CH_12 = 10000'h6d3baf1e6079e22811710f54471ea765365d6fb72e00c7144868ef112cdf26df50a500fe43793772568fef1e5fe28285e4f350ecbe503a3547b99fef063df9923043896bf2b435aecfe7e7ca2177f5f55a54b576e6cab541c1cb87aaf5ad36a13cdf787eb42ecca1cfe5cbfbe6b7876e14a65b920b37751cdeacd27d84c7ea67c51be8242907ee2492be389ddccb9e109e9c1faa8f4ada7576fa0aca0dc3c882b4fc8416bf51bc3b0a8a9606bdf56c5008c078e2a2a7680d90a2f6cc3cff1fb4f999fb67431953a8139e8c93aab3be339ddb12b8301b0b068c8836fdf14b7dedf290d92d14562f4e59750ec60a86272a0eefd31debe5940ee62023d55cf8a594ba12bb487977c3b63d034e6658bcf4b4bf24a9b65f70ae49a1019aa16627dec6bdbaf9e4c3bb64fca6d9531a893a031f8b8f2d3c081935ddaca13495de5f07c27daa6e83090f32b1b0ce97af931e5f69b48792690df155cf402ed3001b7bffed00ebfeeaef1ff408c1959e9fe5469e1f2e24e86c5e957a90b2338536193f88237786f4d059aa50cc0304612464a66122e2c0190901fee67fafe112a7569280042565748488fc8fb4dd20a91301a400de1133b381d9fff83fadb3144d45ef6864fda78163ddc10a63c380cae10a7b1c4214fd9e4fab430bfd0bf439a1056b433e5528df0f9236e23f352e4ad7b0821a1388fd3c7ce0d767edd5d41814552219d0e010c7f521faf5796b8e904a19713755b360ebf428bde4c975472c6f889c93b3ecf1d365d010259664f22cc022e820e133a70a100dc88ac3a58a3fafd3e2d3ea0e1b2bc748263501678a90ba73b82044135a9a6d324d0c53cc0413bed9e70402776858c9b9cc48ff5a5f05b8aa031ff1ef1ae45ebf4f08dfb4e748b1f99132defe3f3218da8ac41c5dbd5a716f1349ec773c9e8c6f5c4ca24147e8d71033c5ee8ae55f8ede25f133bbb2191ad8948337dff42ce49473e32ed5b4b52e06cc862176dfc04b77c4bf65ef478f7b6e2f6a7ceceb584c91bb32b430b57483aa173a18cb9f9aca9f0439a60200413b03aa6afa0840eab8cf55178d222fc5014dba9d635313e2a52ed062fe6af978773647a724a87571e841553e14c0d452e1acffbda8ce0d881f130e62f773fed97af2bd6cde6fe53bb072a12bd84af9be8bd6e1a8a0b0625042952d614cea3b8c3608fb952d4156029b951c5a5cc47575bfbb73c6da4799699692731b43e62e347c09da49e36845baaf7ebf4a158249ae6632bb2a005d74ea5b9f19e08184d2130c8b0a173b5adda6114ccd08ebbe51b1f8a4a7741898bf848020eafd3e35822d1092f96733e2304d125356021424bcc194c5d2b47006346d653236aa3f9602a8c04e1c2bc4b82dc7818164145771e82c304fe8d11c7bb632af63c1c2dbe59ac1548c85060f16abc02d623d70fcabecad72bb0071b368e34667d31de8be74793dc5bc7adbd50543ee843d3c38ffabc6d24721acddf4488a10fbd4d6527af59bb33dfc49c4690b5a7d0c425072e6eaa8304f50c512eb895d657160e6b9d30fc051f75a48287c44219e137de5d9de79be42493ce7ae7b99c69084d0865f4c3cabe2bbe4b7849e84507d62c13f5066d4b81861d4cb2c348391309f4a571d37d3a5ca0cffc810b71457d7701dfd16b7796a422e10314e01e9d345077e6ecb6946d32a571846b8c1dcea593942068aeb5a7d97ab3c8cbb2f83378a6d99f5ba6beaab88e9a9be914c55f39e8accffa040de074ff9c197112c0f25;
    localparam CH_13 = 10000'hb17edee21c0499e11c37cd22966142430120a93689de26835f3fd18c88b47f6b9c88dbce673351cffcc43b695a0f9f308093abcd622dddd076e95d3fa8cd497c0908327a6a9c919f2a9dbda426eb511a3cd44500a0b96f2c2bbf4a00b6e6913c05a3a2fe9dc7889319be6e1e7cd0a0cc0164f96d7c82e5d527c29b594309e8f74a052636b8cb07a321bd69b075d20857cbe19d11eb955c101f5a100d20c011c37eb5375face2551f1db309d9bb722079712782f489fa90170aa0debc44737a2d4064724eec03779ce287d9978a2652e54d534fbf840356774fc2d451d874bee062d728ff7d4dbfe5acf75a8ee1964e5b9530ad688806146061cb0ea6fe3abe9376250b368b333b7e9f5b9f208c270d4920eaa5f72aca144746cdcfbf76a76fa4a64d431b86a895fd11e7f8cb9b65e35963b3facec6350f03393e2069004046eb14f7184dace6ad80bb3bb965c2dc7e5d43dc821fcd07c8c0afc7ea81b7ba5ad634c505a98e9f74c3f63fcbcd028fafe4d627bafb16d79195f35a31f13cd2f78dcad11c3d02103cd59752f48c170d7f2c7eb9b94951cd48a59617896186714322a12b71d760d38939e0d82544c45c0d75641c29c0cc031500e10af304d8e00ccc3f99101ebf7d2ea4259760a9e39ec32d02eef92e65c8ba27aa63b14f6cf5fec84593b58b9f3cc0686e67b9c660affa5c90af112fd035fa64f4a97786bc17b588f35873fc64d059d023d2b822ce9e8c1361d2c0a6cdcdfe37b9931067479987aaa11014d8698aa6c7026fb12cd3a90a3f8806c7c6b35dc90c1877e5484e8e4bf9b78126bd04b13cd96a0b2ebd62532c5409f6203cc01a9613960ab5c964e6edbbed3f73e7e7642e5242ebb2a085932d1a7407231dabff2ee6ee89f4d714c8f40ff398fb96d9efa4b2869945468b5f9763a6ce0c0e0c062bece3c126d8cd4b5950960e5ab3d5896e081f314d3c22031d0f9933036fbe2c5ebd0752b2376b81212880ea695dfb613379308d659a080548435c5b64f349d08780e0a463d4d9b244a75e7971abeedad81c8a62da0c6b9324c933315f291eb16985b5dcab1656eaa4b38ecf7b8ac36742f76e7dfff10a89ec864a55de23be714cbab80e7b8af9e857f3974123aabee8679c7a26617f8ed2439c4b428e46051adff1d192c4dbae0b28c6ba45bb2de9b66a46dafb240b32c67961561eb76ad25152c6971bc1e2f8aa724cf8ffcd48023185984085791524904a5fc79da9bc5d58c77061fe816994186409eb61c0aecfae0f627cee56cbe280348436332bd9582cfe869351a979ecb28cfe1d3a56003006b4020ea1ef9c67319622559f3b3250d3d3cd5042a9c51798a9f7b2e2d55265aca8cdba15ade6652c7523a50ed9114d72469ce4a33f64b21d6f6b7f221561211ac363488bdd30453fd3760f323bcc173c2a45a1a78ba6319c6ed67497618cff67b942b24e59837ed4ceb9f03a1d174b10a17b629939c2d554bf1fc299f8709b8573559abe6b3a8a5f171646c44ea6fae271b4544628744bdba98e43b8e45b3e74cb6d4b20160b76bc77bdbe30058aa802a287b5433c90d9ecfbbaa04835b4d4f45af6988a724d905c3f907c62d15af153457da1f56b7cab97fc4e28a5b88d289da30ae5d112d5112ff4fcef657d27f01d682fb30effacedabad14590095f0f75c93dcdb3a2c29edb2c3841abaaefbdf7af95534c67e38d261223f21af93777f76586f4a62c7782d282d563355d48b3b10edec9463cfd5efb539088e2a;
    localparam CH_14 = 10000'h83fcfa39cb394b4df6a609090346e9f401888f0cbde590aac63e105eb6343dd0f8d6ab323b8f42135e797d99f3233b4826c65e51adef9e3cd93beaa152c2e298f9ff2e7aadc4112f77c91817026d2843f78453cab4e963e0c325e2140a55c735a0acec3f9f94c870807860e797d8af1dc668e3e5f23e326ea17589f91fcc51b9bfb6bbb5353e38454ab2b736b7a5f625f45bdc2f430cd7129414d1bb8cbd0608eb3129347e9bc4a92ed1c98dd865941457ecf6e4d7e95f213d1ef88924c954df94cc0daed8e2ced08cdb2e3b386438ffd528cedde9cee54a73fa97198870b9b0a5a9018c095a43a3090605b190897b11ed0c5b985bdc8c080bb82ec5779a74a309c89e9f44ecb241a055bbadd928589f62a22eeed14e09ac1348f99d7236e9b7e648e9323218215dbf9fb4d4940d20e427cfff63ede39a673048230c492bf2485ec8262948df40e187c92ee1eece1c9bf38ab8f6e60cc9ca5a1c60d50a0971b2db4e66a911b9fab06afed28a127ab1d5ab9d97d70ed3abf0e3f0e0b28be0b23778093f40221b32179e8dbc4f69d2435950e587afefe91e9d6c68a9d66c04e90f41668354ba0750517e3f2ac55e65904755bca20e9dc1e9e10d68dd6ddd9ab3a318be0181f430f09308f356f5e3de0151acef8fd7155dc71007a4e14709a9bb1084763d135dd1ac923a28b51d2d59b0e9e69a66495bb5241ad1ba3733dfcd20e4924a69df80d17fc465a2aa6d605ac334bd6ed2765de6373fdd6c34a32bd020988fbf21ce3f0b286af96ea0069c12074ac5a9549584c591c7bf483e36ae99805b7a7cb93135a1c7cbc589ca4a8a9891e7b2da413550936e0e6411238e25a0ca67a71e068a10fa85431d44c622c9611c256b3a5d6e795fb0580fb8a674d5b1d5566c20d0e5ea353f533abb09a1d3b6181a0de237c3fbd753df066e15ca292ad8b580407acd531aed681b2f54b13f9a1e7b26cae3c30ebdf5576f2a9a47d9067f0e420ed32f9f3897b7d10f5822b891e2b06380a0d7c8b29e6a4f817c47df11795bf47aad3d21582c42f55de464516b5d913f61ca08d8b311e9ba97849deb9a22cb9358841bf518f662ac7f7167a4e158236a10eaaac3680082f08bd24907be2a493460531dd015be075fbab77f4a3ec510b9b97642c58eaed86ec33d22500b1b227ce99f7aeb3c5c061db9f03e78570c3dcce2759a0a3f1bfd889bf448a93207643794a96612a102c8bcc93b8c44ea5c18134c7105eef89dcd9ed26ab335a73041e2ab4a6746851a02b82e7d1a3821fdff634f4991ec53b6b5faf7d76779f91e091fea398b0342fe4b59fb51771147ecfbecb57e01d2e3adcac7cca4a9956f4a0afa7a4643c56445406d85c6119460ed74cbe9bc9c80ecfef53d48d6a22100025ddfdfd9802a00fc6fcfa74304a670ebf0c377c3af3678a7c0624d1a5a3181dacfe8925c81855e7d684bc8d553cf0037bedc7d00b6dbcec7dec3abe193cda790bb59ded9fd27852dfc447724d427fa7129a2f47c746146b76048aae672b2ce0b02f21810e30d7b4c8dbce9e5ae427d6417e1d97345272c6ca591cf0117dcd5f2b16a2b02e5a02eab22d28b9d45dc4b8af43c0107c6a09e5993f649bdbdfa62157c931364d7f25a5ddf9d879d8759166b2f126355955de951424c6bd49e0efcb76eff04410174d9b5fa15203ad69e39a6c3b658e8e673de0bb8eb6faf96dd2e2c86d0a1c1848143bc8a384d84abe2d42476a76b18f1fe89a67d4f5293a653d548e2aa05;
    localparam CH_15 = 10000'h7f8d695ba751d1582461e6752cd3260c02ef7a6d8de2ea48eb134eb1517f11635c3a1a5adb04166faaa9a2a0b228f234f9452ae8ba2261833cc2164dea2f90d495e93394777ae6c1a8e7f60efed13afb6cdd7189ba415f73d0a014050ac6979e62f68ac55ab7fa81d123702f0d0a4cedc856cc911efa14c808da645bd8d09ea342a5898d285eba16f96ac8c6c42b2c962d46dc1c65e7f989c162e87290d19a4e10aab095a1bbf25abb5f837901ec4d5549021a4078e2795f2fab4657b634f8e30cb72fae4a3b3740bd031a07e3e7a6e57579ef4174bf5f2c75bdc19d15f5d74ec96827e3f15b6fc3409620873364ae462e9cf61c6365b3bc93da84339ebf9799cee6c50766cd3fd1f56e44df866039df12a9c0e6cb9ad48e1e2175996869f12175cb93e18c956edbb181ba2e412b2258348dfa615b9d80eee0c30f4db72a10917f5d3f1d9ed570e9b8bf2390928b5857418822e6ad65be5063933dff3f9b3f8ced6d842020f175aa82667b0f0f94ec94dc7a4a950adf0baf071caa490bc9007b2d8da6513d8cc0fe677368747fda7c79e159c5ff440783324d52d156d56859820d6daa8fdfae84d53d4beb09b9f043c277158b16077b096f97031c1a5d7940c2d735e226312d089def07f8b46d5d5eaf872da1f5a084078022fc2109840433f555dd4603149762d689635d6f4b1d6d24a48a825986be732894c9bbf9e3d04ff36e73097577da9a437d9aaf59f52ef03025ef65757a97d74d296eac89d3112fa50ca3621a4e1b2ccf35f8fc20cfc521d6050f993b341e2848bec1efb75f8190d5fac3a5948c3a3c8ef4223ac9f327339ba94682b5ca6875711a99d012649d49036f817aeb49fbf349c060cbedda64f0e8b45217b329ab3e3c75a918a22922ed65cbdb1b42f864253eea35a2e0fc690f52578f66b56c1bd31ad05b8c483768329a427aa30ee93dad893c0630aa29e3316dd743845c9123c18400ea80309a6d68378ef3e3c0150f84a3f21fa7d662a8757c48dc2bee28babe1324f7515d226b101c847f33c8fb065dda6efb0665d2b45d2beb11895ddd77194a554bb8a03596a15bc9fa40d4ecea7a772818f441f1d7a94362ebd49959404ee9e615bf3d078f93ec5d1585e2674ba9c029deb6ea8e8cbfad25fbe96c4627e9deeb9e4ec648449c47b15429c5d5546219c8b9268c6327eec261fad6160dc2c63f395b6ac813318740839007c7a755fb06b8c22d7e6bb490190f8c14a3cba006799ed0751f029092361e8beac03397204f0e88e91bf3769aadc936c72d33be6e40f0cbbb1ca617912e809fd928b9b60e58373a11f6af3ff25493b05d6d6931755c407750a7c15ca91442bac06b471bca78c48f2b80f1880718c7d8f26c6bb25a15db37c83ed5ecc5ce589e251f1aae207d1c1f23c5df743cc72e5415b17bb71c60dfc1c46beef540f611d39ab112b0db10ceef23b63f94a2a6b51e696c04c49016da5f45b07248bc44dd89b74bd6b2efd876319943c9ecf12ce3219f210272b16de9a63c75ca70ea6d0d1004b738bf1ef527b428336085e26bbc3cf3f63beadd6d988e4009671aeac928e70dbd0489657b1e363677962318ffec9aff135d5ebb703f0506954dbee3ec8f9d29e16de484ff6425e80e42c2c3c0bf74404c1ee035dea3b9c80a9511978e946a0b32542145e1302002d5354e5cccde5ae95f402a267c2837ce7dd99499e5f90b95cbcd3f9de348c5f64c2d74916ee7bfbdb5f2c714db44c2f00e943b313b63db;
    localparam CH_16 = 10000'ha35deb8708c2adad762d97bee5e36abb501b28064accb6d6327fabb21bfb690129e6419e152cc5125503b9d168da70f2dc7373238a16ee1a22e59efa0a17f8083553b11c23b5da371527a6940298455a2d7404335b17c597d01c5d7a270da87840835bcac88e92753c9d4ccba97e50091d4b6ef0e2c7db717ab751578cda5ff355b74f5354bb9ec274064a027b0587ac664e9038e3f61a70279607ffeb5ca411b956420498337a8e1c2ccc5a1bcadc8192bc55cd8d6d7510655295027acd9c4277a6ef4dbc087d9d5892126e35da7747294d19c7089f6927cc48a6423b7696b98d79b75295e094472fe3df31e1254a4dddf5a3b9fb4e6dcf51d5f30687602370051bf526184086a307fbf2ab76ac06d1848cc72fb275f07c68b3ed33635266f9692128c2e0cd99e82a21ea7a151a260cb7ef34396045691df263c00face42bc9a1346362c14337ae4b379640596c9112530595e6c952a0fa444a8a0a3d90b9135b5c4445d3f41c2e60b884f1555b6dc26e33ddff77dbac722ddeb5d8e5c6a54d6a82f02a98af2f9e6c99e624e2e9b6950a28a04adacc0ba096eab5483681347a07c9cf8be483e54a879b54c14672d8a66e46b133985a72a64e72d526ddcbde22123cf35c900870d5e1803a6db0d4dabb5b39f3f866130c9a944109eb5c9a235ffa99fb915e515695293a1a2c7da1a02abe4cd637c8a2cedb43cc8f7bdaff7ab64a2ec467b7a810d1685e2cdebc1eb3067615b454349ccc6ddf042985e1171fdc28bd76568cacb3e4d0dd459be772b4866e966e2b292cf813556fe00aa11faba4f842f36ff5073fef7fd0485af37fff9bd156bfc343703f6e31bf61225280ef32a779d05ff43267f8cf9bb7e9474a29ec218e673886ff10b7cea78e7e536daa817124c6856a56e042f143e3a3c00a67c7e2d7d9745893808ccbd8898387d52133b9177002f2514d9b767d6943c9cc8a6c325f0bbbaa92a21170ea1c9f53e9214f9708a6cb6a4e3229561a9a11f2ccd4557bcd447b1957535efab3624c3841f5e42086cc55a1c38dd93e14a039ca0349c82b6a1c1d301202dbf38db9b8a3b67e824e2374696235bac232f6d680c6946df6aab3458e659de9235f7f5b908641e1d2e0d693d373fbf3425f66dccbf362433ceaa2c5756b826f5bff6d5b6a336e968305b6ab747d85eb28835624f2bf7c97db64ef986b2a345d6fc6d84f65726ebfcf05a832aab349f145771ecb8568ea05af9919d252a971359c277b9866d262ab05989c398ec19003ee5f5dbfba9b101e85202a457af6c2fe88f1b99a92c692639c532b93e2c38a0fd90d6e7141ca87e434247e8c6abd8f5049daec472d4d91e3538aa75f35e8914320cec78f7a2c12fea56493dec37f84be81a234f41d7c1a022f27f8762af048b8c910ebf2cea93d6abcfc354c44451066fadbab0d97479b840f3524fb612457b4b79d25c11ab93aa1e449db7e7a2599f03ce4cb3e945d3a0006fcaaa304589092183313318761ddc2d1c6451a04505c0fcad640182c9f1758c88c9381150ac453f08c33b16aff26bbbe72403a67a1565a076f57efef51259eff1e72f54cc650d5362ca986d019fe53dfcf4283513e15e48411e992b9b8a99ba79202c447f77f90cf2a979f3a17bb8977e834e29b87e33e615b7f26905a416038bc8ad74c7fa250cb64b9d42688871740119972936073d158e2b77ff65fc5f62bbefd8d9f6e36bf90503a7bdf63d81604aed00d60b8caad9508429ab18cdd1fcf02e3;

    // LBP params
    localparam NUM_LBP = 64; // 6-bit patterns, 2**6 = 64
    localparam LBP_0 = 10000'h7ae01f579434e068d7a2013010e55f7b2af27d576d96a7947bf0e82a0e87212372cd021a81ac23b4bd51766c414060dad2d253ddd661365dc37febca41b79626cd30f2ef66fe1fb186c8a4ded2f132225e8b582a4f58878fa0fdce6a0e345936c5e7c103573acaa875d72aac98a16d6efe8b7c42d8b97eaad28c46fc773b28e75af50a3fba6823154c51196c50074cd1947e38b34ad47d501960e4b42884f33ddb8d7365dc8818aacfdca73a725d42aa04a85b9da8ccf23c227b252be0eee001a7b8449a0c05bb1773d58c2fba3fc1993ab6be780a83d786972f04fa482b6d0d422fe3ea38ba1d889270437f446b191cb81c01afda706bbd2a4c2634f34a1ce50454b6bdb0f793ad3355be2b789e34240c4293138cea20f0333605bff3034aebe838d6ee7e57986881c1d5109442ddf3e80bdccc29382c4ad44c5880c24d24660ede469798e6c433ed69d2d3b81a1d2867afe09739c038436d98c536635b0667eb8c88dcb782c59b7c19829e1936ae2853547a774477306e6ff9c5ec2e15f26c0a22ebf6ea805b63f12280e24fbf490faa1be2a1f077bef98a21833898eafd3f09ece56efd330abbcee93bdea7329545b81d0ed39031b2a8e1a0bae0e5a362d0494677c046fa952d365517f87c9acf8eac298f6b32476015fba11d929a04e9fd9c009eaf41723b78dc154ace642d7d605cab92afb83d1730e9e5a509391cc59c52b9be5212879a185305b8f65c5679afef9d9ee92df5e9d0244235542350a8dee07b3246bb8f347e893dd7cf2f050de03bc7bab448d052565ff92a5cd210136a6cf8e75a247eae7d80fa55ae4995eb94fbd98f29469a7c96866af57e8c67dd65f8d61277f36a06038b6a4e70846c9ef4d545739ec392f5d38adb00b1ce41d97e20af2faeccb0fd59d14c010eeee75949650f1ff1db2e87e1326494795a0ed8f409def72fc81b6867a921a7937e1ba400e8b3b1dbaafa1c7c0880c49018686c20948278f8293e621251e91adfdf5272716ebcb1f513f6106c7ff930d4e223da129e86c91ab4c6f28cd9972c288bf2014dda6390fbcfe6e7ef77489fd80cdc94a329f917287485dbc347f15b375ce203c4c0498f2474ad38a750e6d291bb5320e840db2dd4bf7b012591495a10da8762822c9d15b94bad8ad646ef5d40fb13732b39ebae2f239f3a760d62ef0a84ed7ed06c22db00448f8d3399532e009717827c3e5cc8fab260838cb34662e0cec83179ebf1aadc2bf384a00a45995bb00f0b2e7184eae65c781e7cbaeebff86e577c95c57db03cf8e752eeb5c2d69b1406d386a6bb5023f25a4ade7a5c84360b4522e727cf9fe8965c613b02f5c3a3b98c8ce4cd46d4a4f4c661d1c202efec2369e922e400f56e87ff864f3f78b9109c12ff200d6000a76b99852eec5827d31d6c85e9059c07dedcf649c81962af648fbfd3ef80ded5ad0be9f149cfe18015e671d721e051a1cc9baa65dfb5b3b887c4e00cc3b37488520f206252f910229fb673e38ec79651320b8f0b7f3c0806936c9938c6654bec402d4dbf778526a53d4eefbc3f9320a1344b46040dc9b5a4dd5b28fce3769f19c0af3ced2d53c53ae8d930917b4738c7f7cb5fca5b6d60b23e943bb3554adb876431524edfcf60a8ff7069d4861801245da9c31ccb9368e9d2b3b31ee5c5fe70bbc445cefbb88737cef338d50918e4a98eb4c99d49e1e3372de2b9053088ca699b059e956a321591fa0bdc1e831f2d4bcbd4691c8f853e7cd09e5e60cc7d46;
    localparam LBP_1 = 10000'hdf85353673c7220df94821646cc02db267e59d77d53116a54d3085d52a0bec75df2659c392a00d09392c5fcb47a70769767f0b076d67fc3370659bf9ea4e9a17484a63e152c7b66585cdda33d44ea897cad4bb1bc5d9d6a69914ab2e4afb4fe8c8408e2b501d43748bdab4ca382a96db2c7348a598d2ed7e6d2a4f81a6a00c0164de371c146d5b57a66ca1acf91346a16eb27e9dcdf773548da4e1862679e2a47dec0f551a650ca4013e635325ffa9d4bd4174d86185e7792798962fa33af30baad4791e533cc1e0dc39cd9c199244e8ed3d1c5a8370eac5b14f8f76ae48eaa89523fbc7a3424127fd2d69bba868c54fabad48d9ba8d61ff09d59d5c5e8555f2572928680318117d63595275c3e1fd296af58d600dfe2da9ca44738acbd0f60440a70277c48c826a706252e48b6177def3d3aa19602a094fac1f0a4d40f23efa30309fed81999f949ef62b7fccf109673a9dae9ed32645777223c06d8d9a0b69d373a421fd8575e6a425cb8dfd034e68a15f889ba3a0b81d791467604ee44c40597ffbcf55ea074cfc1d3bf26cd6be716514ad44607ae9ddf4f8abd718f1bbe4b5420972840391b4b093df3de4b819bf0d2f8a6364cec371649b6a16d029924d7ba59e53653753ad0fb6f26818c1ad4b6f69a0d2ac731a24ad608b8a581213d73b2bc5d8ebd4c2ea36ad04d40211533f536e29222c4267826aa6e724663f764ebbb8ad65157ea41d30953514dcdeaf2611d9b0f2cf8b4297f3a1975d3716b90d11de2876dd632a53cbd6bb46d80cc408be7c48710499af5a0b00e60ee73ee6dd7b93b02de42641d95da81209148a7659df34ee9bc1a9a1519c56cd1cd9cdd3c6b6481c7ed91596d34b1f558e3a1f59ae58b0877d9554d68002b14958948c1d309dabafda07ae50e66388cfd828d67a70df7c9d81ad78d84f891463e09c853841b93c9e2f7332ec8b3ad1d3733d9615f14167e47cc3337f66ac2696a323cc52589b3b918c5298dd34d8efa88d7770f59fdab4c6184356123f230fc8d5e29ccb0dead7e4ebd01ee89681dbb4589893ea7d7f5530f09043a092771188fc9454699df41ac014a91afd21ea6fe22f11b172f481ad6b5d4527ee15cc3a50cdc200bb7c68b98581601640eb2f47ca681d35d60d5588ec747dedc391a9d1fe9e2d18f94364ae560eeb61ed3bdf89d4237ab8f3d7252cce8d56eedfbf6c41345d6cbcdd4ceb6fd95efd0297a24077ecb4644607a93f63c22c7613961b371362697f2614dbd5ead429e67a7b25784d9050c7616a43f01549a778ec6a4191fc9aaf7b8499a42995fb62df2a29dd655aa0232a20ea09f6ae8bcce487bb8626c1f2708c022567d8b785da01361c548d966ea18ca0649f2e5a2826fe5ffa304ed26a42c96ea1294a3de1967b2ff2aa5d931aad75c5a426a5c3a337d0020d7b07f8ba9dec2d05074ca39aa3a071b683f5ca6ad3334f0d5385ff3d5774323e210ae1c17dbdf2241b989279f2ae76ec048877d3dfe3c6857e110e38c9ddc70d1363359b50d35d856e8a472ef6adbd29da7c892381878c93cfaeb414cf4f0f4002adf2a697c86af947684e3859d4327ec5f6bc88d3884b02488e66abfbcb312dc97bfe82e86090289bcd7337369f982425cb4f4f1dbb2806422ce8b8415c6a20ce245eb4ba6974c2c34e57bc6a7dca04b00472da583220428266fc0d177bcdeb25b27fe3ed92f0212d1e3ccad3272a48087436616141b78a9e9f217fcb9652da1ea0bfb14a0025e76f49ae;
    localparam LBP_2 = 10000'h627c4ea4a60e5edabcf1e1c61f4efa08d5f1767fa640131cf1c6444c8e864004dd20082fa0caebf52d1d1f2da03d77a45e54dc4173b282ab6fceb02bfc1be04ee4974a57f90fbe62aa30a0e312d8a61b31a4cf2a3a4dc228da2e25ec7af77cfd5cdd4c8d9d70edc0a1c3818e0e165da0ac7383131918d077acd27b3271827be865aadb9d4b4360428104855926ce4f29b564f87ade57f9ba6e0aa717409d4276f462466055bc3adce27e216c55ca4bd4cb10313f5f7d1cd81cc4f04e34ed718f7e9815f5232adedcf7d9d904af766803e0dfb80b08e6b9a2f33bbc4889586b3472472b71e6edbabec374869af99b1d06aed897ad12b90489d699e511905caf4150c9af78741a55e85b7745fbac015b8244d945f9bfefb2bec16976c643c48f70f68aa547bf74526e2cce4cd6624255544e60f7fe50bebf9ff9cbe6b20411b72f863c43ce6dc8238b3d9980ed4a5607d0491a10c8fce7bd04c703277f870fdc89f3cdda24d4ee85fad405c795cdb9652d406a5c6e3f33d04cc0c4430baa530bc4908d5a6db5f4dda4879eb5c8b6eb00391c2238e8dc22b88450abe0a2aa96da9dfd85fe2fe79b27a2eb6fd1c7a1dc1c705ebe52d964fdcc2990f4cd2a8369267f32ea024733df2212a3d3b2bffbe8d48634a915c2f2a5294ffec2473feff97dd425a7ac8cd6f4fe2c812f9ab57c1ff2e2c1d6cc3b7e2a8fa32e574354d85dcbd185bd35e6eecf3a3e86a5cb992e88ae95beb5d6ebaae2a428bef7e35875ed70c3283244fbc1e6afa044616f68594b59a56d047e440210f2bff74bbed234c1358337ac5136b2d0c0f6472436aaac7cf086e965a1d47aff3b4582193133528a17bb70032873def423081d145a1a083ff94831fedc3a0a1fd287c0467dac9648967616055adfcb68f1cf2fc3fd6098030bfbc4e2e0bae199547c633287488c7b1c4d5b0326584833bb75f4d891cfefd7d5c293377fa697a495f68fcaf677ac037b90198182a29b6859545c84923f0f3ae9f24ebddb214a61b57c60f9cb390dabeb5dac76890e60c64332b1290dd08f23e8750cdc072b758ec9333280bad0c0e5fe426fd92b71ebd3a2822f0b56bec7c2bd8b885366344f02330a9e82c4a9ae00ec37f66a30b624e8ae3d44b3718d3da0b0d706555277d7dee10c8db4998812182988b85669f47dc413d9c5a5ac57f38a32a60b0d5b9f6be72df39930d2caff154ffb149f860cca2cdad5bdc5c83478faa486fc05fcb948f2eb220e0f8151b15591c6443f86a66c645f22d5f3375064ec5bedf5afa6b643bcc936dc030d000be768a937b88ba73230611da2e207a695bc4518fc8f6b444fc44ee50d4d9cd18caa842acca62b947544b5a57c8e5cdca857658af550e8e6cea13a3ec4ba2c02ba3a0e5940c3124a09460b9d7800301ada3c6de457240c2480f89a10ae1e2199a97bcc16f110bdbe5ec84b51a3889a805339ea8c180f8d697485f954de591a11ddbbc12fc82922cf25a35df6614c051c253bd22853eaebf535ff44c79835ccf041a6a9c6a56ad0ea83c41386db5e28df97c7022fb23dfa9da3c4545eef470f6931cd082a1a35c2bf25a882e9db3437c6164356e1821f3f696246da1bf6b4507598f3e2345d778123fddb9daff2d03976757e640873b2b16c23d2233699234f5f2f98cd43c28197dc090bab6cc54d4c0cb0194e0616ec7363abec3efd1907cbf98de86a85ef320777b54be326a249a06467a8f733b7722c26273a53862d006993866fe706c4e;
    localparam LBP_3 = 10000'h71e6344a0856a9aed5a31409617ac943ed9681f32fa7280d464debdb89fc40e5887239d1ad94fbbea68168eab624fbe27edcd5cad4d17551f099d16a3ad02140cabcea5ce1f622af471d82a3f20ddbaa5457f2fa78f5b7f233d989840446cc1dbd9698c382385819ed0563334eaf58f3447b29ffc30259faee29302b68c858d58890eb9b040abe1b8fa4024fbbc8f0613010edc9c82a166d5bbb84d9aa482ab4b5f155723e289b277818e7787da187ec2cab738c976f976bf9db737f5c597474b21b7daa9a7555edc476850bf38bdc714a86ea006c51438ee36b9a28a2374ee62d299dc4654ac8f9febc026e3a24c99fb8433a8fd6e8a47b8bddf9b7a0322350a179a8ee02e8502ea6566d9c30c2caff1b2fb27c5775ac62e7802404821289c0aac60e54c5106a1ad63c795b1cbd908e31b94c69a901cc742232670dba75f58bdd1edabfc1c804454faf9020aad60a280c8c95dd88ce3cc59c98daf8907316b640621b460158f3ebb00df254b9e61dc760f89333052d2c1bb061b8519e894205ed4e7490b4338657f801d1dfbe9fe6e25b55b2203868244f11f8ca5db5fd17deda0c9d1e124c9e45fb45bd745bf7df42a462f470de9ce98a13bbbcebbb6adad6c76ad6cafdbfb7573725214832c340fad8fe4a9dc86643c9df6abc6742d48495779c297cf2e4a9661e3db8f9bebbfb9b18022e4a744bfea99a8b7465f07d87dec4f008da25d28fdc8f5368234d3b5082c94b144659b81747184038d8d1581b60ac146b41385bc2d25c758b56ac5e64ba350487b3c740c5061435603f413fb997c3690525ffb6a4318093824997399dce438ac22e8f849207a8ab7b050bbb1344630597dbed9eff1919e723d27fd483b6c7a9a3ccec8d2ebae32b60bdae152e850be50dd2f791fe17cf9980dd6509fbda1035bf47595ed9de52c07a0179f39185e7008cecedf5df7959bc7c89e7b9f202cdfadd0ecd4224287f410440e8b90c329e6031d1f4aee7af54cbd10b6de386c5cd6032fd64b836c9fee6d8a0691b9050d67475edcb3ff9f1f4ba6dfc743612bda38132eb7bbc0acd114cc1fa2baedcbcde4f8bc665428864de5bd4857462f0dbab88b93ebc6aefe0f301ad7d9ba6090fd5f55c7ea9dc55677b45e3653d2ec05d40b32e760ecbf549b140cd41d6156837e194bbaa76cc5d27bce56a5a8b25a666a1ec0942f1235ca0ef764838cdfc75f19d00debf0b70e2ff6cdafb9069914ea240fcc1dc4f36aeb2d5e59e6f6ada77481ef8dc16a4653b0e501e5fd515858a2da976b350159e9bb2f2a935dd4056142e85704392be2c4bdbe67b871105739e85a873ac4212781d9006d428576d735db0ed92c95547d5dcb3e4e31327571491353e0b8ba97244874f5d7eaa7c13e7c4a68835d5e491c96a5ec66ab72a41dd8a1d11598a69d45012e01fdc645e06e9b70698933d7c50bc165299d1a82f02e227a6db2013ec2dc222c8c17fa9ca4314067fd65cb1e1e297646a0e113e6ee968c7ba0b353167c297db1430a3d6eedac37f5897a32bfdce239c91fd9df542451e01bd332a16680ef74c313b2338dd4217027ef230eb38cbdf781e26909f4979a5f4756df231a1b3a21da4a56d40729c36d7e53ad541aeceabaff1504b648c235b6a8e755c511930eceb254aa00e91c35138154a2aa69573963402f823c8200dd023f75446f4b1a6de543fc5ebb05166654392950026c43e29165e2ec1bcd3e496cdec3e49f799b82d4b0a5f04d210c9b89c865632;
    localparam LBP_4 = 10000'h4ad6ee94b1820cce255bbce7afd94049af5c45ed5d43dedd0044bfe8c147cf7d22413b5f1189683dddcffff6c15f8d2dec2f0717a02e858b377a01b14e7018340aad3c4322ff580ceac07c708bad26022c5b87ad7ff791f5033435d0f011e4b568e9c34d93f54b42d962dad1dc6ceec2f7163eb84e49ebb174d01db29061b389a51b68f669031edd716bd178bbfbdf3cac4f89ad0f75605fb337d70073c4785eab09c51f66ff8bb939a27d6e7ac02934c165ea66c61aa55578059ce64ad6f83514a3124a2d7f1f87a10cd0de29711d2f695e7ce4e92e3adc0593bde98f05f651f2f3267532104131dc0ef52f976031c60d0446bc03c008cbf68b24ef77dc8a1bf7af5278eb502bf4fa38da025b84dd0d6726e877c9db6ed55692ad949846453e7872a1fdec051d21b3557d69a75cea6f0fe289dc53110c0be4dbcfefde016271fb64e69d2e58b1a9d38932f7720ae5b598a7f7deb494334753504f932b618da6a4dc16fdbc9dadcf402471815cd8e0ad5f608937c10aac016cdd10fe91fe27d80f12641086459871f49431cdd79a3ccc40bea82283cb8a3e5c538dc249e2029d8fab5f08ee8cedc6c45063b5c70bda64e0615afaa7a0d93d67aac61d470c50cf0c059ba35625a36566b993504892770943c7819092ad7c9b154f80d3f828351cd6064b85b528ae30f591b9cc3e679b3e4fa5429bc4a0c0fafaad003db23149ba0ee6b86d8419dd87fee779570ac6fab8f2e71bac738e1e915e141544e95a6b556dc382c2ed4a1d894a3f7aee2d8d67d3465aa3a19fe25c4376bb93a652c54d2aae9f7221065e052f2461e57107ea9fd09cad624bd9604fd04291c43a585520a36112500b217feb5c8580676061ebc09b610ce0377f43b661f09cb97114091f2a9def4d1beab903ba8ed7d1fe03b5e49c7ab7264e9836526c8abeb9400acc73547f71823c4bef5c4d6ee994746fac703a7f42c94b47bd63c0aaef662acd9d5639c81b6dee853af495909c56885ff00cb7be70a74af658099d41bba7d5688a92adc759850714a98ce38a684bb4522e6bd5538fb1a55817769c59ca362a57c466f1431ca5563f0b2bad95bf6ad87765fcea2b5a604726bad6c7bacfc6815f5d2326857b3d7ce2eda029d815829475c732cc189875fbe0aa1d9ec2385198ce1fb27a8f84edcdfc511a89145fe4e685c140c283c4183ddc3d177b6378be6508824c2726dd1a340c69b109ec5de840c305342bd4a70ed0d38455d6e5e6fb992dc44c16238ef679bbbd962ed8950f3e1f76d8c33916fc97ed9721d20260c7108a4f4e3b1e1d86baed8b0a64c5899102fe800639a45570c686553657e4c267ecc08592f65700b0bd44db2cbd7c0bc50a03bccaa293e9514ae96c750f9ba69ece4c3f91da0b76c2e2198015a2fcf413b09cb9ea7a87d6ada2579fdff9d409f984f10af9d7244b653577128cf228c319e223a08bec31ef4de98802b4edc28574b4a2a914ad718fc934f1e5d6e4af90ef38a377b55209dbe0464d7ebb689a582b61d9e159bb9c25cfc63ae0b1e5ebb404bfb505c8db8f8f39f5740921249e62593773483e17484d886b1e6a0ed51b2275601c411dc9d634f0b71fd0165d13e93ab36092fc86a956da0ac8083f41993a5c32d0b11634dfb963c6c0331ef6e96d6c0a07e612bb258f637634862d7dbc258f6cddb1a27f2b81bbb915d85324d9f3c8c2ca6e95b0dff6c5b7d1b253017d838434a1a09fb1b3e8b984da32e8d8b77f25abc6042986db78;
    localparam LBP_5 = 10000'h555fdc79c7b33ec94c616b8ec273b440aee381bc45f6d672bea8daeb408758c0fd0314ef838e3bbb880e8971055bc1a33d96411c509959a52ee20a6fd11aea6ad0a49de4c8406f36391efdfe1a22a6b2d200bfaf1f20989224bf019d61953835835885fcd02c5a2619f2bf2a35097ba0b013c9be3c7b3b9109dddb12ca61e19951dd94e5356df59aa3b588fa984f52ace655ac4aa6b87e4377c78841d9abf2e7a1e29759fadc7b2acff58c6d4cd1e5bbaf2dfedab7af077efb1ea30882146ce8672a273e654de4265fce16e228f5cd622fbac101212f7f7787e4d50441eb016b2b368d347ccc7dd54210819723b17762d230749f38fcb2083ade12e5a24220531acb01fc90d5d09252c504da19c1417197416d19d2a1fd0c3307cf41abc271908ff0d387f542ff289a816a0f8aff140f2721c2358f722a6bca026f2889f35295a6c3fb26cfe8d22b23642edbdf850a15966c1e14b75aa3bc7dd1274b82d665ff0423d776e4e5099a07e9c75f911e03dde25cd2a35e69c011fc9799bec670117f925ba9dadf0e3e5a1f021f01e4b85fcd187c9b62b1ecc5a1878c658ed5ce5d4798dfd9f9bf21facc3eba74de8fcada6932661de499f5997d485d75bb9d5294d64d5af3a059f65c44d57680530f661f0d8af89bc37671a59e02fb5db78462c7e5fcc4269be43799438a9a2b33914923a328f8a14dc8cdeecbaa807562fe3f5124dc576715aa3f16817bdf01ef44672a2f785fa80c4bd82919d4af2a4a3d1ac1c44000b80cfe1b1ecd12835f752d066ecb8f360f0fd0304d72da8e8a32bf9d8c4df2686f8ee635f6adce9fc21a99a296df57d5915fddb47a340e44c3557fd968987b4197bfdb2fe006818ee3e002a80c22928e172a64e87c3bbf04139969ed55e789449fee6f626f94c98f7881b2222021be578145c3d410075518d282ae6f08304ea8c9e343494636551f29c5ba4cb1f74aa70b216f5cb7fa6e61a8427da05509f5b2dc7ed2702f381e315dcc2661c865efeba5916cd768e9a0b1636434979f19544fd81d9321b3ea754178cf79d42252593d587e30b499f683e2514efc1f339d4453d24dc612a813421878388b1c4d51575a6c13cb92ed4ba725b3ddd3fcd2ccabc22faf55cc75d4c7e9190536a56abc5b53247a457b42ac7ca1f4d6a7c3d11bcbfaa84a384b858eb1296109dbc3c00c0a5a77fb60a9de428f1426828cd4efe43713f6ec753a4383f1c72f6f909f203466761ddb9a05d3ccf8db4664cb56952e6d8a3975569652f5f21eafe5b99b03e1bf77c983f703492ef9a3e37c615227e13a19a0fd0dd0f5d33f5bd0289727a69a9427e068f18c7dcacbbfa1c2542299dc132d2441fd843a73b14287768979854c1172a62236be7ff358772557420d8f0dbcfab381bc46e2a97ff565d4472257b0a28c14b792b07a45c3a8198ac052aeac52fe9fa2158fe25b830d51eba5c90e6d071b0a820ed3dd53a65fc27d0ae148108911d49475e1659e0d499f437ab31436aa213d1744b925a2471543fb8a99d1a6e49df4b0d75c3f7ae17688bc0a03a194593e96a8e361939aae8da8331f015fa6521a81f7226bae6f57c6d18b0b709cdb09280486ac9687bd127831c5c93ae0b698dba4e42e5b3d3f839aa3326b6aec4221124249ba113d6dafee45a9a0d12c708ad9aefb6c89abc86ddfca6a556b56d5c49d96afbbd6980d552654ba0107f5e7104e80e09b62a72419fccb8cca5787ab681e4c6842521e179e5b621305b7922f7cd8;
    localparam LBP_6 = 10000'h3ccc7c5e2fb3524ad780da83e830888936aef7687d615a642ccf1c858b2e3b92d6ad62509c8b07cfd2522177cad9219fb49c24ba9e913800681605070fcaf5c4c10207058ecbbc7502dfde204c8e9901d86a92b7a1ce9ec3e711ed24c3ce9e20e805579bb411bf63c7a23bfd14068bb23ab7c1907b4e1ee9d033eb9aa148cc20821de4a6fbeef048775c9629855a3ec30cf3b74630f21c4280d980384d47166c91b9dfd4a0fbb273ce12acdb33cd1c5349373dc339ada2088d91a9f5e31d3066ce7a6f6806b688c24703f72602215e6f7168bb66dfa078048e1a83fabd9efaeef02c22b213d0b7763b09bfa200dcb768892ff6b676e64bf89180458e83f9a864abc2fe11611a3f995f1f9db597da5aa3754a9d601d6dbbf3555cbab6adab5417abc8fc3d1e808b1ba59594d66afc643cb287214f6a170e87398280d211d783d1ad54e6ffba61fe85c3372f3bec78158537be51ae69d35d105a1a628576f426eeb8069950a2db5ee636c819ec4345be30818720e5484b5b8f87dc9bf4b36c5f225b25817e439cf3a589c4894d08c66fd291a96a13fc75a9bf2ee9df4b4e4b3d55fe2c544b9f907f309676874c2fc9f8022aa8565218d7d4f2483c692a283aea9272367860007788a79454a7044da9a23dd1c42c00a3edb3c8d56aa7cfacade9be000723fee3510ee78f33cba2c74511b72a295de3867dbf293004c90eca61b658b508bc0f0fff73ae2c362c948af03fc77050b250c5cdb96385b99603e70a0285cac80ad41be77176ed15f52aecad121db4041fc5541a5f88348095bb40dff89a7dae5f3fedf865d9fd3b36528783297ced921fb87dd7fa60d40fb6c829b3c5081a262b7f31f21e9ea6ca3846cc05b9b6f43153070eda3af305518ed674dde3717f12f62c397dc4571eb266e8c6468269b7d9c9268dc212a432ef3f2223eec077398d4ec5c0b30c2f74d7c907d48acac9c7f95b8a72ed7a7cc931b7492252072d1e110d33cd1043e7e3d9a864a61f7dd493dd0a026bcb6681183deace8361f87fd490e794e792bbed04095c6ba1ae242e1ca4b419301f86c832751832ba6101f3dda77008f5ef3101f79300fdd4a3bbf2bfcaa0aff5fda29a876b886be5fedcf9ab42b602083bf6df3fee3a6b5430c6c3fb9c47b8cec2c5443baf271a37c072ec767b8f145bf52844e6c1fced3e9913e14fd4e1004ec4015758d7604e94e361217ada453fcc188c648af1d1e4e2bd1f2c5dc0a840110681ac7b4afdb542e6100f86bce724e2abf46d4cb635ae302e1f9a7c449ecf6935813780770272ae0373e6efa702307ba536afffa625b7da0cf1f06bf2c949ace88d33a6181776f499209634f5f8ca6a8a841e9a311cce5bf71e97cc7617e334b90de5872574c3aeac920924b9d8d5a59d1cac0e92f9b01da0e5f5aad1892db3e6739ca1a34ad7c1b4c1dae25762ae26f8d039ea7c65bd4583f82565828ce2682c2614fcabc659a46a41c4ac8ca18e2871b045033e290abd50ef2ab7c9a35b64c455e7caae715d7fccb80d8553c05a9b6cfe1f1d6b4f9a19870796e1cad1a04c5ebfab177bec722d7a8d2bcaa181cd98553775cc65f921884ab81ec57f50283a5258b6e986e2ab142f7da6c7b828ba547abc15d502b369446c368821741b9f9a3479a8c174ff2a7c38d1c9415661f0be1fec3bb78dbabaadf074ae4a5b57117fb8611bd984e7237c5a362557b01a99a4ea45343595377932d57e549d2c11c5a66833aae623e7160da9326f6f1e;
    localparam LBP_7 = 10000'h168ead0bb6e4e80451be70f1a3bf3358bba6155cd1c25a586f72d751eae046721fd8d34e665d4131c68a3c779f49962b40b6eaa6006f37c982ecf01cfe207f6f5b3cbf273ebd81f2176f026312c384c0a04723366fb1c52303aa962b4b997a0836e3b365a4b8fdca932ca564e40692b1325748873cdfe9c331ce09b5ace6b499bca97d7a962ad061981e2a2580a49a5f1df6d2097f9756017dc564ba7cafe1922462508d210a130cfc5cffd6922ddd4808fda3a0002cbc2ee674ee61896eba3854bf9963b7f55815766520d0167f6a4c343074937bcd4eed9a9d73549ba189e7485a6890ffb93a73acab15fe498499f315d170a7bb6eaf91c1461e55d7b8fdf5a90bc9acd6a82a82d86da6a4d3fdfe3b22d50a07872570bfa558977e686c142d37210d06e2f92e5dd869d799cbf1a2b0dcca411c8e203164e761809e9011f10534d551c77573933ecc9d55a16a51f4d1fadd5cfeda5a2f69dab11714eb17922668a971a966a63d29567b0fc23dd3d28724fcb438f760b1dfdba788c051726e7186aad934b1e89d3a41519e41fc3b845ef06d73536476152fcbd2e27ac5a595c581939c2a2e6c0dc2fe5416fb7cd6e76b2325e86b9014116bcb64001367e47a5eee1a6ead8cc93d9a507c462e490abd526a5c5608bf5b452cd240621c9560fded25c1727356b5341a1d534e8f37d1612c65216181aecea6f90ebfccd9ce79553ece0f3de6331561275f92b92df43306bd3f6d8faae89ed795149d891982143ee6de663ff41906203236f7520d79d59f5fbc2657448e347607616cf162cf7a70aded0c35e966ba67c428cfc0d755257db0708c24084184c29ad9a89dba733a18da8ddcdec2c32974bfbcdf0b99a7915cc1f626bbf7828dcbcfe61579c48902f93bf095f9c04d3fa6708b9c82405dffcd82ed9f6dd5566330c3362609f02999ea2360abbb109cc094e4fbeed26b9e123495e624bc5afc3ee9c67ba46df7ff8fab30b7fb04479fdba539039b08d6619b7b01b8210b274164f6c326833ee5b803f51464a809128fb1ef2eb438769576122c445cab3de67cf07e2c281b4c1140f1407c54d6be4a9e234ed663aef73323d69d47d1c2a228eb5d93954829589a79aa441925810fe8f1f98b0f1fe0b3029bc43e0f41709edd502e35d182961023212ae24c71556c566144e3383b7efa23595ac8b77ba96f2dc01f78be7f84fcbb44b44a4bc59a7f6099b2c87b2cbc17b11ee73b8ac2a9f0a99134e7fd7c46e3d60a19bed8da221122e9390b9bc98fc1a87a6645a574701cd77144185d52598483ad4190a2e2406141b3eb3bb3320b65c4a40c08267b2269994e37859c060547de0694f39017ff5b4e326534ddf5a36b9ddb887c1d7c5e0d4ba2b041009979510233732610200f11f04b7e2a456e77cb1cc8f40cded062817b9e723e6b652df07202fe9dae931c1f9f5b3e587ea3c08a399e5f3377a61e56c217ad1b63e08eefd89f713a13bdce9a074b91bcd92ce25facc398a40b517406a953e22cf39bbbd26337c2c451fa6e869f8b35b2f288d5a8ed66c1f3762cb75383f837a54913f44bce24a9f58e8d15d1236f1f147ba68d7be56d31e9019bf8061495db9be49a1a862335814fd5d15c51f6f039f0f8cb48c80daf93c992048658016748a0e7992139a704862284c4fdf6031ae415b39ccfbdeaf7e89ae62532128cb69d7035742ce74059569356bd3693ef683b5dcac8e1ce7d0df63ab7aa9c51424ca02dc695f487dea10ee7e9238a;
    localparam LBP_8 = 10000'h3c3a44c28081ba886f1873facc24ddcd907a6cd7096c283c23c48c6545285aed6e1a894f1f79b42b0d9955e63d8e4273aad6b39adba37dc16d5a1d6b8776d8959b7294f7fa4ecc04641419e9fc6529652eef00adcab68985773efb034df8ece3d78666fd426a9d88872faa715cfa456b436f3318b5858b32c4660fda47bffb1e176723ce8ab2a27bf28f61d0e1994ed489294bf67917e65b291d7ccc28d1922d270452d3045a72d3f125d017df1fdcb86f689b9a220cbff7c2e9d4ed0915194d4af95723c6ce8f5c53ace61cb9b65411c34f34a780cc477a3b72e3c027535674af8969bed927b83ee23c60e2e2fc20a011e84e3f65661b431d522a573667cb929086353cafba380d5f51b947a007adee03e8f5ff334b320f9e9dedd04dad9e359820e39461ddcf3cf33ee585922c164dac155a2c6be8c11fbc8a18b9144a48cb28a49fa86d76d3c485e5b2e5d63c2c2a55e0cc1ade0000d1592a71e20ebdd1cf3a90ed07c37e76f26033727e311beb485be5c39df07338f1b5a8fbe2d4c82df0473b472b7f0085beacab68e7b5c696e2d52c06d1caa44d6692fb866e5d6af8fe5be6ef4ea2dc2601d830d33dc39a0a99f6aff52f92da27f2dc13f81501139eef27b266966db63407901c20f8453e3334f044668e4c0fc197f36a6be8f60e2bf4bbca96b0c2784cb357b03e7d967326df4ebd982140402e9e2aa6bb8eaca57d4511295bf08b70719e2a342f0577ccd04da5bfb94f850257b8654fec49288c3bd84563dec0f1a62f2f97f188191b960f6a1a90f58861beee23c945ed1d1fda026b19c01a96e578e44769d7b309997f9ea431d572e674fbbf9f3d69bb76877d2922fe5209a04fce65c62b259a161136b66ae470c1030e649bde951d06800fa1a3f0ca6e5dd1779359d7555942440a831958012d10911636f072b1035605207b40ab2dcd15a85f830771bd81983032d9c0227300e8e240d2973bdf093b523621db9001253b24b3cb66f4822cdd843a145f265ec47a8b0297f86ed932351777c245c1f4ae8ae5f13416e3231680ce070303395cc3e33818a777c2c5a11c6dc7bcb5471c5c2f765bfd538ceeb6a9652f7896d2b6348abde479eae477a38487797d95602a1bfc84223233ad48edb28e8fb3d2e42bf78b53ac96a7e1ef26bca9094ba0240f3ec02106efce3f79263781dea096c08c4fa78a8c8127e6103844f956950014791a9b3e956d5cae85a0fbbd694bb348ed28b9ba984b66467c4629ae5a37927e3daaa03286b9af7074b4ebf331c9f5208d0b6e0f54e5560fa4dd0502656bda0c7f18485e5a6c253929d9f43302e0232547db1f210537397c9b998206889dbd657743ee55f6158597f7ecc28b0675bcfdbaa31e842efcfa419582a43b2c1cb01dd79036459695707f4fb4eff5244187efd4ea5c673edb2adf87bd11af0c7a23f17022332bff8ace0b811d2f19e8fd9cb1e451f1922c996beb4b2665924b294ad2319d9761d3e20553dae68ef3749bfe924b03840cd4f87d834bdd1e041a36076d16885b95f0d6a3d71001469212199244f118c01c64b9efa2fa3127af28871a9ec4c387f9a6947d49e712f5f8513b43abe5c7db9b84da67d2f2110637d9b9ba63e1bbff74d96302700d1d5266892df54977734ec8cd7e6fc496adfb135e00cd2ca24f16b03ea402638aaa3d137b98604cc9d703b6d7b58b2bf68d71b633276043fce03d13e4f99bd2ff5b509f14e11c3e13629c81a1fe2b9329fbe112c296ac424f6;
    localparam LBP_9 = 10000'hc53f18afce5156a3781dc74f4c260a7b9b232df2c499be767cea59194bc39ee22e5cb07bd7dd7e20fe0e5c22508e5e27b572724b8faf82bea5a891ffcaf53b2f50bdce9c69cf9b296540988002aa805a6c1965fe2bcc10587630dfff769fac97ba44989c1f58942562c82c829309f71fe5a606a568f814a21c13bdc9eb70bd588bbf99f5f53b38fad901d8fcfde848211aca2356a2c21184a43831321f9e26f59c40f96ccc48b7922c70122298570fcc81e9f03db0f83441517d475a669a44ed5fc8f9c4841f3a6fba44222c065c79007e751b6f36e7a624bf64c7f7661021cd923f6920abb1b29d076c4cb18168c55a0df51abe4ed9c9c8654421984e8ef33349b6051b6811663ed6886474ac556902e3f21ec3bfba1e6df486ffe87cd3dcc5dd5439df056bc7a9030dab0b55dbf245644d97fdef9bafd082c29770ea1ffdb8538a3af3d6163f5c08e0c6cbbad2bf22c7f6eb7f95b98a3ad068649782b06b80dce5c21b5657dab706a74c82424617cf8df90c824beab3a98dc821bf449074954a1e5622ff4bb86e92d48836497b9cbb46501e4af694ec3b0abfb7caf71ee4ead13913dce1d80befe9447dc21a6f2093cd40a4f506d33c8f698d7576db9f301ebb15a986a8426267d9307e6e6fb055366a47859a22e4b742760156eb700c6838319185edc2e59354bd75ad4ca5741b8ab5e6247066c9ce7c311ef43aa7087d326a7c6e9d2ea0b1479f2d8cb10c592cc1c354f4f3b7fd28671f3133694a091363e3a04639652020fb24eb3973b9adf58ccb3a2f49e3f879cb05a9f2a90dfddec0a8c5d9e84d9ea175cfccae5b698abe3c5ad6edd530d42ba618ee9836bbc19af2c8b6c4dbba8e1777081c72906dc04a43c51a64c326515441453362d1577ea0b8f765bfd28b581aebcbbb1d4c52f8b02fd696f4434878745517007f34ddf05a4b08b73f34001d5473e1518021c159f5b9fcf19835988ff67883ea767e993eb05a7a7f1c3c11feca6ca6781f0541810f4ac80115f999b66215a2c352d54780ac223ca1da83903ad39b24f9c621ffd6c91250b6e0048b0a4a422cd53d28f5d40cea81099bbcbce987bcb746052b462f07bb33d79646e0d1bd7e4d0870c1b4d3ac30e341f3535f24f3ebebdbfd1c69b09b704116c666d51efda0baf0101112354bd4aa5e955219e583a53c9451c6921a0e571de91f5f826ca42d2f352989f59b72a6c2f6599f7b284afa024142e853c0ee390617d26884dfdbae707e7d6851c57c18d14233bf1aa61c034ad83044ae58da5d988df9bc422082b114678f4311faea066ae39796c839a9bfb3acee63c8fce084096f07e74fb2711d482ced3ecf238cf3c04d38df5ef53c1df8300fede4522912c0a23c04543b6cd9de0c0774f31c0eec253178a5ddb7655c36e89e3478fa655ea5660e7557b65cf8f9e5cf7c55ea9cfbafc0b6726c924638d857b350d0f2d19c19a4c9417d83fdc6e73898e44dbf29a2b30a392e6f782e394d88fb312113449a6691bec450fc67763c94a12028c41e6dffdd1602cdf6b7487edbe2682a011045de615c3f1e8daa7a8686c6c1aea8ddb68d79655e263390075f597c0b1f8c6eb0bd0c21795d86d4a40dd920a2bd7bd78a4e40b1f5c22e3c44b8fe37d01b9b2ea35565af70f8723689e6c4e34ffaeea9838a1f96441e439b48e3f86c9ef09ad5a42f9861b684dd58d699b9c42ef7e04222fc1215a5fb764c4315c35725973eb4ea079b5b706902e4c0ff24368462f38293176f;
    localparam LBP_10 = 10000'h3de4cfdf54d8d8833de2346aa8bd467016f288390075a6a06a22277da5e92d10e31d137a8242137f49eb448a60785c223cb636af08dceff8a2d2fdc5d5be455c0245bb6ac6c637e63c8a95b26dd82c0794fa67478266d549dce2ac6803de83ce83ca51163c4862cf177d8ad03f869a7608c02855e2722c63a7f22cc59edaad82ca4f644c4b90a96d3c644b89cf451000629cf5080e72173433b438ec08baf87904c455724e11f939bf5850d3b1569cde9a9d9990f1537c7b18243889bdedb08bd0ad49a7656d5df0288cd629936791fa9d37f05f93ffb26b3f16b067780dc163fde01d171019e99eb841fee5a25fc3dd5f5bf93b5725964ce03af530f8ef8d03d3e110d7929ca65474505d294e97fdf4b105cd03cb1c5a3edce7dfef41963403e94c3c02a3c6e616000ec6b55f9abb323dcf5e1dfb0b70ac69fff06aa72df026bb00d6931ddd2a0703abd6af6c82b5fef9d7a7564f769f0098b84302e0ca6bcb47e0c5f16305e18876c5b94175e91305c737d6bfc0d47262981aaa964c22ea72ff2edef2cb494286baf01235debbfd070f3ac7695eebeb96283a072dea379940ad3844d9b3f135ff841b8f218c69361b5d276092bd59943ef9e3b7db98c283b1755db2f36d89bc02a5e9d43544b839a04e6dfda1a27444e807d5b7d69a252ea01aae1b41be9215d0e3057ad9b2cea9b6d1dae19ec96700cfe15b2681193aa8e4a3e29fccdbb09a03bec805e97e7d1561f5a6829c44ae58834a83197f8462d054bd52b9ddd8aa38c0f57ec4c7345d0ac53805c19d46abaad5672696a4448dbd60a7fa6ebe2ea570160fc77f234558a27533855b0927edaedd88be97ece147e16aa2b72634499b8c44a70c9f5053b2e3837e54e2d2deff4e0ebe8dc8330577196c4d5aa928a5ed51e4f4e355aae85563939c1cdf10ad8da022cc611a0d5c27db21adba472b97153b718441846ddd0b537fadacd4d2cfaab24a0a43c0d9a528eed66d965ec58308510f782954534a48121d882879bb542415069745b207a8cb67e3f27d14144090c57e88782d44f8924ec8de4d374166b5005aae87b8ff6631c608ce4a3e2983a91979873ddbda4e554cbe70162b60275832b3f4f563b2fa66bcaac8cdfbfabe74fab609f2f283b6e3f49964722eda68d1b9533562e595cd0c76aaa466c5577cc56d3ba52a37fa20ae134fc601f981ad093b80e15f939cebe062cfbbe53002bd6f486043b8ac3ee44f9f575149874990d6290923492d2d2c804373541abe5201fecc02e1b1c2059dbd6f9ed0c1bdeaac00dfb726f19f4e4d831ac8447ac9e1794538288377dfdd1b23902e8043a01d96327283329ff45067b9a6caa01e4ee7c0bb8611b49b7910e1b95c5d243391b88c957e0ef3c6cad9c5ff3157cabaa3d1a873797c5aebf68280794aaaa85142bf40ded43b64c796888e3d85b66a6f7b87fba5218afe6de49cf312adc936b0209ee01633b58a61b335e2a393386e40994052d15ece3aaf267ef23a88bb22a2d7212f2df7eda36c91de624716718d3762dff698f2cebf86e50c1b9eed518909e6d532e9d9fc93393db895a05ed630663001b438bb14bffaa6066da564ba6cf47325bc203bed38d8f8e0098ab3e42951469df0006da83a0e3a766740a965dc7eaf6a740a3e0eaf38f6fb73630f79aebadf5ac1277b300366da4254324fd2ca07f114e70e453df9cc02b08789064173737f37f1e8333516347b283b1db8f9b1a5a4144bbe6723b9289d22d8756cbb4e8f;
    localparam LBP_11 = 10000'ha9b09568361c917678317f3c53fdaaf8b661254f3f49a8f9d7d9cdbb26a4f90f06cb84114f7b16e96dd1f01e6690a7fa6f29cae5501376252941facfc86bec1641efc3fe29b008aafaf2aeeb26fedb04ef0768cea91d7290da3b5a716e0cb291fa29bb1f422f6d261c5f7ce7d71f04cc5d91a70a340c14444b9b4baa3b0b0930474dc0415b993cece4275df0225be5c44550e1dee8a8c91fea5e128ba58153e7008d4ee4f04002e98d09ca990c9d2a1959ca45e47f76dcece328d60c62cf8a2b62d540cd2274e5e54e8d65d996556bfb95d56118bc11c375d720736806313d98198f235d9ca7238a57432f587078f11c51097be01510a057cc6a9b9592020d3659d47f8c93559e00f9470df0aa95e31f95a5d02a68048231438350b0bcb0392f0c02aea3e0bb42b67827170d2df7f3771c64a4205b3d59b454f4497ea4e72b2b9e26b161ec6df5febb9e703ddf2797e686e642f5966a90e62c17f10bbd57388807fc506feb3201ac969517f73452aa5122e6a66800263377d5f79168e8d0676638f3aba528a850eb6f44cdf5c84bf406eb125e99ab3d17382800ca4a08cda34b9c578737b1a2e85457137c967b7c5ad9f58e47fbef6419129bae5e4be41d741c7a525d767dded61db9275554653202789a946d1dc10f97414cab3ba0c629366d708512a30159050154b363867f815f07f885a9d6945812306867c917fd86d6e91f20dbc6a392f7f6f747dfc0cdeefdd6222c03054a464cd1a0f105009b1205552d572b5868547c2d28595442f8a26a581fb22dd2751f0d41e81ba3c9bad4ddbf40cd9516954240edc1466fe32c74ce44130f8c5b2eb8e556fceb5bf618ae57b256ea1c3d3cf594781b5b9685a9f4c6375d05fefeed7e02223ff6d996db39c5899d7beac7561202540068df2c86237f7e6a55413ef63d9fd59760ad5806c5fea25536de05fc089528ff35029ea241cfc8f53bfbeffb96dbe41b407a3bfb12e00ae3d7c797098071b216ef242c14722c85e46bf82b262f084f1e3a034cd6a30bab2c459b62432975ef18fe44a29d7edcae3c5a822c33c94d247c7c97f3d9b67cc7c4b9011c45299064bd4707dc0f23ff2506b9d31fbac53018179baeb9eae2801820c256d20f7af74d20ebde8397368332457b6fd5f5d7b3d29b4a318c7fad9b9d7df0040746cfc0db959df0b0e2e8d3901bdd1bcaa8919630ac32b01c115274adb4fe2b6e52f9d0f90c5981e0a47529b0810fcf8b75153d9380778a8493e287c9175852418da89a9292c7c3642303a4f7fae6d6d5180cd8ed2bd0e657c3d1d94f49b31dd333e169952f8e32d7b5b11e0340675c8474fa35285d692bffff76181f25264f657fad7941f117102f40e0c8d3123285c0e2c4e36cdb9de37455d01c67f75eb265abf0471af106cad02102250b6324d3bc25be79882f42f07dcf50aaecf480ffcb8f4d262649dcb92d6a86e219279ba1256fd6e63866458fe7d2205f71353bd40f07a35ebd917070360b3e511559af6e435c898a474e57112dfc67da2bdf0ba282bd818e486ab973e08c073455819bc1f51fbbff874d74b82b4f4cf957faf6fd3efe173230acc8f10a7d39bc8fdc1a73f409c9b122025671a81d62efa6603a5741e5295d52f4abc6dfe753fe155d299af1437b1dce53d20d2a3f637209e01f8f0536c9ff77707ba12f174c0fde4b585cd2c907a404128ccddc907373f1f916749efb5f47361d02c721a0606e0e7c27481b091f42ff534e1c9b95dd1b0498ad;
    localparam LBP_12 = 10000'hfd56cc5dc780210dcb7ea05268a0fc06d143af1244bbf203ea1bb54b073f05b9af693740421e7abd33316564855751889964eaafc0dfc7ebdd5bda6ed949a3e306248c99471464e84f83c66af41465968783382ac05e2fa4066ee95c1890b67ff70b735ba70783aa7007353c21fd2bb2131b254213558a42ce6bcf3875b892f73a3797ef17258dc29b7da665263db04b93c554cf886f1d9f2eb22469c90bb818cb7fec1d12c2e72aba1510f1b886648df0792dc84be92a3bfbf60df10a298189618bf4e4337542f58723e47cc69fb2a24c2f744742dad979641244729b7e71016b306bc949c352851d29b44190c97e25fa15f9475c62b9b4397842994278e4b7b9c4d3ee7e2bd5e59113a7eaeef02f5251e3251e4ebc37dc9fab20f5dab0e9aeadbff5161aaa997d457cd60b969f60d9f71e11c67dfc09d33979fa31451bf31c93f83884b84e432820a4ab075d06401e3331439c2dbb78b87544b4de6c1546ff433b746e9824154a602a73ca763b61bb465f1fd917bf099ebd089e4eaa2945311ca390e63d54027a99ed077180df2805c140a4c37f366b0839c26d131195ff95ef33d719a3ab22c8fa52e933b56301dc0a31e835c4253fe3d9b70e5fc1b36bf6ac965bf4d412c95a53756655cf8076cb0246c68c5f0bd31502f47e071f101c740c87ca4e5f376876242bedd18064b9c9dd6339b7dc3ca30aaf9ca313dd263e2c3eb1bfe01603c941953214f508cfcc7fbf7af78f81639b5c0da6a36f7cc51d6731b60565fcdeb0157877199cd1b847e1b1a358de8b26876b58eea8007adbf075c79df8e5a20f43d8081c230da33493754831736ef58dc77fe9e15ccdbf7668ba731e26ef0b9cf132a4d67d4e8c2c97eed6ffdf1508801712f90fe9e5f444c4c75e65bde403d5570d2428dfd0e2ac02bf01e005870203b1120b558cba4fff4d091605ebd5ca698e0077bce548b8c7ecc44b9c6e2cf8435e1046ad6415c54666e320b0a9aaba17d8bbee1ea19fc1b18f4a35dd0603293a34b81391a2c8022c61553abad4e9833fe4d341b9ec2847357f2efbd0261f8d467bd8490afed667721b9899713e4af1a81026771a4a8a58e9ad57fccc83859e7819b8dc8960e8419746ce711ffebad4ef138f7a24fb46d7ad34e1caf7593e80d79edc5188e48b502e45e2ab544744ec83cfa3e1cdddb0170779d04a21c978c9d7cf357f15c9ef1d1c5694640b9ed299fcc027e67df415154c3cec5bdc5ff9410429019ca6264130210b4812cdc1d176778eee91524ad1e1d00b99f3ad67e8ffa0766a673338fa1450396c07952a2c368474d12d6c471c98f05f16328db32e46a69196ff09cae11f18846ec95fe23842bd5818d544d90750ac06d2b0e36a60bef2fa539594f7c003869e3c8bfe63dff5f301526007b3ddc71f628149c8b2a179c3f6bb8ffd37cf8dd23c2589437eab428800aabd8c22196c2af552cc55961fd5a88f52197f87c5cdc58b0997414ec2bb41dad30f72b9055a00b441152c728a357b4231a12fa0198dcdd3d8dd3a7b4ed2cff6a2b797be95882cdf10558c3c7968d31183f4a999f97f1f2daab2ea26f04c965b37a99db541d42d24b703e45655b645ac098de7e05af301ecd3744a39be8426332c805f5a0e7c828948916151aae1fc04e1ef93de74b64e2fbe782d996a4bfe0fade72727a02a66b0fa83771e7faf6a45adf2ff831cfee5a65f6c072d0ce6ba96319690a21670aa1a27e4b842ea1ff060aeae5154a8e157736c883d;
    localparam LBP_13 = 10000'h3f60b4bf88650b7e89349ba88b326aff9ae0095f457e7d9489f59282590f6e80aa88b8e45f84b05dd02fe9e1319d1160e3b74cc4889637094677064b7ed3b52620bcebdfbc76e3fdb2b5784282d6158dcf87b493c868d048e09ac4beffb25526bedd5add6165d2f1adb9c7b36c757e3db85d7e4fda2f50afea8dc1e9e372aa303df94e5645bf805ec2abecf59f17b2e25c60b858fb12fffd6bab2c66b9c800d9b0bb4b84246a5d82fae55c0af133027d8fa6fe133a76243495de11f4d66c287b7c41f53ba7c86327f4f80e02ccd8d72efcf4057449980bcd62dbd6ce6ea9acb3986d345381128c92872c26268ce48cb0e8bc80524cded545c302096c89f430bfcada17a3993b06c6ee4762af48fca9c3186b8db59716349d89e3eaada163e63eaa0ec11ea1749c3d074cdc721d88719367068916b5ddd6da0df6a252e5c7771a12027d46a2fa96642b4f8a043d4bab1321f292cd76e799e94abf8a15e5fbc5f1ac7bffc6c736e1de0c67beb8f4b64a3590bf8e98907d678cf4a5305c0139b5074f0a8c35e5d19b6c533d502a7ed20a8fb6269d55f5a6b2c589f737bac484e2134a2034ed60b3c20e961d87f867369423785c26408225621514eefb9aadf71b833403c905e44f7795011fa14c6fe821ad4dc9b9e1334ba9b5fa6bd347f312dae7e80ea2bf9ee5f2acb4a7b5763580b5b635571345b0469f7c8ed8ca20da50befa60d350bdce5742fb7103e7a647e7921b5dc61b97f74312ad558f063e685e4df699e86add5d82a9f072b96ea1ad151007948890e2ee58f7b7d9af7568db8d978faa142f050487d335fda226ba8767e3b4aed252df69f5b0daee5c7105c65e1c19b6670a95d95a537f0807c5050499c40df08052378b1491106913dd74bb172d3c19432a08bf7ae4994c37efbded2af885b3164947a3f8ee74d48eacd25175504828d3b2f20cb5f867f98676de18c5f2631dc0e1816d405c6fed9bc77b0d822fdb2b276d2f2db924135a8bb22c8256235a76a36a8329295a4d16fe1028fcda6a17bfb0084447101c955b3bd1f6c03a8339186719f35046b68d3179041bf1a97a3f09ca1d7f76e8b8e47b9405583343a36f7678e59679065bfc4ce56fe6d168bfbdd2d35fc22c79d6956139e7bab73291264051e71cfac857aee50faac034a5fa298a930ecc26d40ab5b88afdd06dfa030c2e74b94ddf1e68ec6468b40388365c3c6d948175fef2b29ccceb04a090503ae5cf8a48d4ffe26eb84e860790cb75336b53f749bbbc365612bb8cb2a1583c11e0012e908438990f84a2a818d02eda2a5f228a53e3ab40157502a9e477b074e4123b38800dba6a81c89e9ebddcd7fa1fe793e642e38f8c28e5acc39313f7a2abe2a129cd69353154fee8cf4f11bc3db58695227ab4793646647f3d4a615987fd45c1f68ad7d31a1e09a38b7f22fa730d058166a06615a1eaf1086e21bba958e21cb5194a6e55f0fc155fc7d5ca12e1a3bb652bc06dde47c60beb84f9d77836898e7aa7aa893a8199e2d3f463dd06b1ce6a22de595c486b67230afcfeefb31e54364b3b50d4dd2075d095965aef7354ea114a322d122b0e3df74008c0f060209690c4c63c4c41106423be163d9a3c30f0984703fd0e3a662f17fd2bbf00572e203417666ca586ab0b2396b70682e61a41d4c04c8d3f4dc7c1733e6050a46025178165b08defaaf85ae760d3f44880198dcc604bb7e752ac1800405c3481b5957793cee7ce49b889af9bf8a9a5471c5895ebb72b;
    localparam LBP_14 = 10000'hc7e0f6673d8c4c87c2ed03d532bcbeae9d710c6526985459266b71ea32ab830a1d10f48d9b2ff70996af02889d7040c6601ff831f4088cba0f5acc66e29d5e51a7882be0c5207ec8b5c3b7bd1bc6adb4e4d84b102f8601cefdc716516301c49364eae4b942802fd767a61c22beb5ef136dc36faa79a1cb66a7829aebb34ea4de4f09c010e144f0d17d7b77e69d59afa6eddac8e4e5f592132f58d3e004a65154e0903bef45d04d53ee01a1abf806c3e49c2fbacdb7a5f45b548ac3e617b6afe75d8c4ef43b4e9452e0a5a0aeee39c3b96a5c845b6d60e3abd4b751424c58b3adaf4e384db295282cb73fdb5b4c2bca0269937cef3980de1b8190b0db5f0d73d2ffa20e03c3e109a313b12864c4a7345fb14e61a90bd4fcda70016322dc0e41dbe9e85709bf91f1e6d050e7455f21122f17b80ce8ed9c97d70d902ceba255db039fea08660e2fc8b10dcf479dc19bf8de77c5a0bc2c58979f7426c3b8b8c6420c80aeb768f38cf6475b84561a7d221dc8577f5d761c7b741e5ec9252a7cf3851132adcd299fafe57743d2279dab58d31c925f946df9ee5588ae41b855a3bd2c3e8ca7e9f6be471c1ad291c1f62fecc509dc305de9c4572373183eafa9306788ad9769e37850698691c1271d35fd4768960f2ba50c739d82723930b02b09f68b6187b7c02bd335004624826512d930403816a9d9cabc5c9469d15cb2ffa465cef13f13b49998fd136377eda17272f6be9eee9d3eb27720ac3331757a6c9a6b7709a6274ded255e3a848282f3b2cd22acc9d69763c55a2d1667ad9f2c9ba3f82879f3fe40af50850c950a4795d668ed02e842d85bc3a6591234a5342426399517dc694e21687be2bdf4eeb0ea2da3125367ff8cefb3dd3932c98c31702b0603d695dbb9333a86bdc70ecf636d1f22d4a9bc47c557bb2dcab3159aed729e386be926cae373855155dde2c66a988ea5a9cd40d4de3c521785a44dbcc3bc6251273399809c21bb893ab6f8779e866b5b5b15c62cc57b04a7bb6c0f1d8caebf9674626c42ae2298b3837fcfdc9de96a15951aca55f1f455477e90df30672a1b87d0da828c0dfd2a0aa6917c1eb9b04755117ca76de61932049ab19890d6192e78acd219217a6a54630e43c25d653a25e8b7a9a6384cced96d055996d36f8aeb0accf87c74678cb242db263100ac34cde521023c6eb73e97d9b98191e7e8a25474025d95adbbc53eca8035ee025252b401f63c43fe960b9c2f80aa9b6f6dceee87fe42011f07ed491de11009a3ecb93762c32da022fb62d8740480ca57d99a67b6771ebe306c6245b20988558f613e509497b9b047fc69dcb4c11bba9f01a95ebc3b3f603b57a288586d67b1295384a7008174a9e78e94fbbfa20722531a76b0a46608f35fc7f0fd7632be00027fc7c649a9244e4aee1b9f2747a8eda8c710bd225350ff22617eb3c9676035a05c7394dc94153ea9a3b122672edf2f13bea4c6e925dd1f5702d76c76ad336e74541469ea9942ce5eac3cb515f8df0962e2a1cd175791cc58401ce7f228886cf6e0db05631f26a985b49eb3a89f2414866b013bff3e05b1528d73969215c54dc92f1e395d96cb7089c3fd46fdeff288fbd9ba74ad545c4fb307242111901adaa9dae644dd1043258eb478578c25f0c71ce048fda9b83f9bc068f2e83c7cc477f20d54374b965f2fca80acd505941408fb2fe86239509b41b781ee0a4e542f5b13ad232d931f7b670c16ac3c78cb0ab7d54b6ab4e42c425d24e2;
    localparam LBP_15 = 10000'hdd669ab788515f39af77219f383810423feb18946c8dc815794d16f3e8027e5d9410f313f876a47180415b846600299585f6768bd48a79969942a420fda78df7788aa16090ac99b6583e60beb7bbd808c6475b671b3a63a398dde24379b3c83cb8e4b0632f35e8e84d7a6c45ae6547a75a9ec09bb261a5654de8c7cc9cd2fb881b08e0f44f80da9ac7141c7501a749edf988da1855eae2a0c8e817e02836ff6d2eac0ef8c1487d8b3332c8d9bf358b7ff445e024774770940ee5d8988201928ed913dc8910616e38aa3d14f2c7b3bf33c15b0c13bd3a37c0a1b2720adf145e64172898dea57fab0659c7694fc0bc7b3c039f78958318a0d145c3ac2d3f8e431a1b5097e0c58eeb78a49c8bb164fde5b88eb5c3630125dc814a8b6522f86cf79521188dbf7609b133f0de28ca650d72ccb1c9cb3a25c8ee1d14d4235a9097f54d62979a82301761db79e66093a631c8be32db02fc98ab7a58954989877aa6dc51e02db9dd246ccaa7017eb2cc078d7f75d3c0c92aeee450cf60d80b9724095bc62cd2100afcb8c858b88c99ba27f84ead52f326997bc57d4c3f35fce6fbe29c84a97b7a3130c299542007e9d3cba9d2cd8a929d78b00bc87a6b30722ce1b6a7ea7e0a5c046763cf7c6386ad2d6752976a8d16fab116f950811961ba7694b725b9db5de57a237fc9e45ceba3ede7f411319d7d93919a1b2c0984874f352b9868b09cc2f33c2acb94dd21babfdb9e7794a01ce56c39abdcc864c3f6b17b93eb9427d0bcf3193c4cb16835e40451fde688ad75afae5490d455e3fa2306c7541361646ca6e514b9ab7dff3bb15eab1f530ccd58d6b229c6fafb2c7d98383db4392f4f4651b1ce4c472f46a9471a01ba177a95396aabc9bf793a28447ae84f5d7eb0ec9550f37e5124d9e93333e899314312900d359f6dce6a80d269aa9ceb9f7cc2f904b4e84e9dd8f620cd970a11f89322bb4ab7c00b922a3840bf45b8d7d62e6042fc527e2a329f8957db002920651e34bbf23a943dc87438830f210aa495e439f86084f4c8fc9adb8f535447dfcdde31b95128112d4b74484ebc3ebf0a6dc19e1711ddd4b532b6cbeb225120eabc6965e411e4ceaf73275565797895f659d8c75c7d73082b9109cefceb79c18f37b60ebccf5944ac182a8172c7429c7b364b3c5a3627920be41ede32ddbe109ac8a4820c3a299abdc8864fa56e2ec4ae2552c019bbcd50e8a8f7c07ebe5d4055d700bf42ee73a4eb9c2afa9f3f16c3ff7cb70114a99c7e675d6bf6de5e5e2ccaec1443712c844cf5a1b153ab36eb9de190bcbf5385876dd3709e24bf9d1a2d23f8284f741a42e60c2581f2a3f24adb33b2308d4cbb5a8205c97a552b433c307090f9a180e5f84a970d33cefda5eca3d65fc46cd6b57757b3b2ed154b24c32c5bfaf5f926088fdeb29988b7548fe6b8f598ac4e35d2a4df5b39f72b225f7ccfd447832d3c202e14552ecae642873133437310d37684b25e2c8f48eaa9830e6e7ab3487b34d3936caddde1a72f6e2e0cd268dc45377f7558cdf7590f4a5b0f0cb6f31faa3c4f4c426f04d99c6d268eb47bcc21297e36224f73dcf5af12f425efe11ce02b7070491fd94b78fb698e1bb651ae7eb9b90dc81348cc10cbe4c5ee01e48e24480e9ff743043be625c4e23ae36eef41902171242344e2c1f9f4c6b7745b1a281c18ac8940a8fc5f09dac17a734ec800368be6b70304be3226e655725c4ec28249efd127bbec02a4bccc119d35556f0f065364f0;
    localparam LBP_16 = 10000'h4eab5b1873d902130d57b65d0e9f8e9d8c16ff4551d60096e4a8d370ed97ccc2b23b555402b2ea43da12a77790f63fac18ede0faa54b08b8da327ee915a1ec60a00d5bb07a4353468e6123359a6e51ec88f2576c48b1b5e5cbfd994847c032a213c0d44e8ac16cab89b23a1e015ff59f40b7d74efcf76787f53436bfd68f3d85a37267b59feddd0300ae7a741dd3a1170d76acfee3d4f69001b877618c963097a25083cd4c61a33d673f9c74363633676b620bbd3c3495a9302c584688efc50fce786de63a359eefe3d5d8d777b2813e34999e4ac40143cd73ec0fc4e0b9b82116f06d01b54c016ca998907263a13f98ee4cf56522d4ee8465847e18aeefc68117edef080ca6a4b7e7e06898e70cf84911a37226d5a7be0848c7b132f46ffc87eeade99ced0b624d24aff17c84014c3745e2c2d55e45e1284b6602ae3271cd41517422babe74c55dc60a925485a9ca197c76d41a6e5395a3b371d5b5c230807384091d981eced3c9e72b07a48f1ecef518b07ee939c4dea8fef808e808742164bddcf800999b985bf0a1019756df4ddf47109c1083c3ef6cac46666830c8aca9aac0efdae713886d8da00701243ab59bf48cdff898f2443c687bdfe3f743c86f42f77d5b2d9acc7cac3d7f8d66eff0e730d787ea8926eb155e4fbbbcd9246a0804448e1c08d0c267be410b5845ee7294113ea18c553fd12b34d4532094d56d94b8581f3b48f08eabb5af2eb99466064e247dfef613acb9771b34b38fb0225bc2dca09f76ce684fb80967c13391b3b05951a767ae0b44276df37ce184797974c7e4aea6086d4dd52714bd4914154696d5e2c170becd926a151f01d0204611ecb4a4e0077f1563175fc097360d84e34286737b13d5dcd10c6b8d05fd9acd91d56f39002ba61b3cb625d86ad1ef166ac0157af7d32523ed24eeec709a5822683a12281e640942cb48cb3f9e087f42280b5adde806170484f935e9541ac3f74010dce741f331e841e78ec14811f97ea78349748d3a562973f2121bb6ed3c4a0bc7207af0925d67e22b4a61361ff40b5cc770c71fb3941114fdc4910f4286d333cb83aebe40283d559b80369fafa688fee7fb92f6f76524597040c01f27892b0448ef23aa4cdbd94c0a8ad26a644842b8f742972ec3da4b7b2f274017687f9467b9b268bbab4bfb1b0086da03005f9577d92d86fd78758aecaf1a0e581906f8d49f27c582c8496f1f32d5025ef90248bf643fd2cc6fef6640ca97dff86edee2ef948d068dd70c9bd496e7181cf4712adc22dbc2aaad055436c3ec4eed7b33bc042d55463c9f609dd139540efc6e08ef9504408e08cfa0bb2f12df28a6e72ba6633ae9b0473728de169b8c46bb3a26dcf3e84f0baf27fd52fa9f5f35ab029003f7c396217672feefcab60f9b8ad09219d522d7a166ce2d46ad5b1772b9ce233362a4c4fc1c0d86e8d620098ad4f172b3e7128e06376362a8699c34a0706476aba85fbcb3c8a53f8589c6198baf0bcd76e0f0e14043d04015fc244487e7cc5285dc99eb8e12c9f9cef9c55921d15435c6d2945dd7ffe3d77fdbbe927b46c611275d464ec3e71b2be8072fc086142e8abfd85f623b8a1603e2735c0ec6b8335c4368f0dfcfa02f49f30a81fd761376d8b58b5d2fd33c8b82619caf4f3597e6e6dee2b3a90e23241a4f6e55fe7dfe1fcf4bef4f18340d84a153cae534124b667b0502b6d9932433c4d3d8fac37347619227365def6d5a1ce197a6efc57b9b24645f5ab776d123;
    localparam LBP_17 = 10000'h2fb52d12db3916e40ddd0b179e04d3b14197abd8a17201a69be74ef671ffcb26ab76c999d0c4476d6a3320a847ea66034e050d805944c806e39fc04706f1b1fdd2b44c1ed9e0064d910d56cdef35815178c1751401c8dfc12f4484857671d537558d491b900c52720d47fc49c33cf175e425c787cf3cf2cdace137336a37383b07da1e21312b13d577960afbaac25d17e0ebc058bfcac185a090a801c2298707963210c88b3f300331ec83c662878e87d9f8bba356368cbaa2685f4d5830130643affbdc76d742d9262595b868024cacfc9cb4c8c99fee4520bdcc2e04f67c8d53b4da11b60c9eba5fb8d0d56ddbf25c06fa2d3314b6cfb7e483d715c6606636c22f00440d6706eaaf6b2917d440da5506fe66794bb94abe639613bef39794f5bdd8dbc8980e84212766a0f943d2152c758d8766428643e5cdadff2891c29333bafcd5d2c575d4d6d8cbdd920739bd4580b9e69649101cda0be23edb39b9a534461d078ec8bccceaf1334861a8bd4a2c809b511a5888b7ef389454a3c8580486a120bc5069cbc23ee141f76be1c35488adb0903e3ccb834975eafb6baf50e1ce9f3fa898ce189d916dfffb3c63263afd7c2c71132edc791acdf3c325cc86bfadbc29e9b305640414047119f1e014f591ed8a99f6c3fabb36ead6e9bf50abf0cf6de6207b8d38ac2648f03f5d5acf6d79ddf8c1acc3ce5f5b057d3f565c73ade6c845dc07541c89aea71912eeef575d63aac99b510852382ce96222ac9d14c73e1f54cfd5db0c5d5cdb79d5fbcedcfe1e4cc75cfaa25b3f142f76c167cdff0326147d0cc3c3ca905b7f5a1b5b2c9e49748f4f205a79cf5a342d87b320e4f6c4b1cd40164da3ddfefb7d5a48041fb261a3a605eb46f0e08867ae9065c61eaec2e650289ef74f053633398ba7e368e27bead5e9a787a17e88b402beb21a77eeb90b9e145a015ae95ff981867c4081b8b43a675a0aed4f51e00da7f1d94b2ba318a437ff63c246c24eca24fbc303996ac806c578e9171a73ce1a5961f418d4361ffbfcbdd57ab8858445e993c22c64d4fb17dc41a85081b19d7ced61561c839ed1974ef12560ce942386dfb9f0b76bcee79a9f27227ed65ed5a284ceb7287dc97e6ced8d8e1c7897dac4a34743e3b7fe92c75de4f8ab8dc145428c9a12a213a8838befefdb41a65731ac24ee93c3fbd6907bfee9b1b55014188a8bde3eb57572d59d6766eb94706b878f77ca95d4ca43e6758a6c7487644cf3863bf7ffea5f69e2720037f560946c66060273227897f400c01414a47c809b4555ff96d362af5d5416fec70d14dcf822b0218e4212c2a06163ca8d07d2ecca8e87e8a293f2750b667f8143aaa4e586acc7f226772b4098467d9151ebde77f913b15eb56aa7547bbc79b74f3e6085b3160ad9a0961e8032d36c3b10e04a7e0fa1ac473e64945e1516da9e73fa95a78ccfa1f889101896e070a69a4499a3cc3a7b7dc5fa80256d6589c04d0b632fafa595b8421a55dd5fe2c991eaf6c9acf3df1e09dd19d6b6cbc272af0c79889779db5ba3ba9b1ae4b2246c4f82545ab377aa5e468d13338a6155722e7980f286ada63ce44c800fa0305e406cdd000185f2d386075cc09cd9d14ab4efd951ca2f2216da0766487b47e28058c5f87f304822ac94097e9ed0da138488c6c1f9af5dd0d47850bab1c399e9608131b7720efad22cc18a21e86965de5588a801d493d0cccccfd128109e46168b4b6853e71944fb73c77e633f80f353c4f3d1e2f4;
    localparam LBP_18 = 10000'he3e48043a52f2b3f7498f1da9af42856cddc8a518e894c626a7e674b2dfc3aa278dde65a0e2291d16b8f809c9aae822470e8f81ce861a7512ff8cdca570ebcda303717b84e131bef73f5ef152a6484180684c30b562dc2d9c4f49551a1bccaffb13cf64d123d8761c5fafd95cf00a5a4631cf5ce665aba00bab66401e247021190c70f1794f293b7fbdf5e3d10cd89e93614e4a8add87b85abe4a02a43c38dd91074497eb3b20a81f924516ed1e5ab275edd6df9de7a3bff0e0d29b0442d799785d358a7126c97fd8de3cc7bfc186c6abfd9a1b9184db4265e383d0d03c898707953c147d9b47290c6744980431d03098713e5c185794ed73c77e11f939cdde13bd4df9a97ecfaade278baeeb8e88d14a58c2ff500bcfe53ee093c7f4483873a73fd1c178b86e4fe08525b349fa640af589b761b6bdb532695b73bf521bf197c6e2efe3a8e07964193785dad6405dd00d822928396d3a96f2e5b1b3d068918206aa8b0d6ba4e841768216f04e4b55e8c2902e9a5d7a59d0bdb1a77d4b05935f54ee75c2ed1fcda2db88d11d59d802fb6b9bd917f58a0a720e8b86c4518ab9611b1c494af4cddecf9b7dafc266b8adbac77aee684664b9d94b21c456626a8d2560937a03756fe6834f5326074983fe44faa9ef0bf2fad3cab43d4bf480172a1ad69097662c1311a110a2f63f8112cc6835961f9cca1a910a12db79cab597555ebc5df4c31d2931583085ed7b60bbbc2eefbba321864b95dd51f9b70640903ddbdf1407e20756d5c4eea4a245b851a6f2fa1f3e7181c46dfc6486e6c0523e7c06419c750aea697b234af35671546a62fb55a794ec98d2083721c318435fc34d058b2eb8aa074a92d0872a446256e7445b1569a8afd847031c073b25157bddd09756ff66e7e68685c4267758887593562c01dd177db143d6269db23e72081cb39d34d287ab99085a65e749923c15c5ee1a3b364e9e82ca1a19144b24ad46dd3f6811d30ed7c5c40b7f791f2529a8ecefded0b42dbe57b63192029eb2753cc1da20a8c7490c34b9849cda75f1c4cb0671903dfae2dcb0178951f75e776075b60feea24e2e319b65add774120619c5e1290221c2ffd1d7a224115eb9fb61f3ad4e75825533b4ed9a4d7c87f640ca6120c23a1688b08fd2084e4f37ba28b823a8ea2f7c77b67052aea3d5f8f85ad5c62455fd63b1dacb017b029f1723297421851d049830f297fc33177841e5ff838254f572266adc61d630850bdfd990a061b6cfd2c924a98539d1b810691e6cf55e9f3bf3cb5bb69569fc119ece7c6abea24931789b66d725a72904beda203d14c39903933a21bd180551d0ab520a09375ee7dc00952f23b8f35360ed5a421903f40f787acfea62b88b6c0bbeeb62dc162a4f113742a1d23b5b0ff80b95df7a0a0a4fdb3c5ee4a6935fd725630296692e97afa363f6343fa44aafb04beb5825d08398db3eb1be0883b3d4247ce0d58325ffa73c67d3100e6c873ecbf7d4e191b4ed965a8e91d455b994f11f1852f0d2ca4f03f67f102eac6a4c7d5742b1fc6dc080f98f7afda28607aa3da24f7b64c523131e608295f6757d06f412a65b8df6f104a325cf989e0aeaec523e2f6adbf212d42560b6fe701c6c2d3088ea3cbbacd75ad6e044bcaa1a1a4d88fed2148eed6f6900112212c492f836145fb8106e19b246c58c6f46be535549e95344de9739c940fdd6f4e9053bbd3461b8a9a240baed6312c6397b93dd492f19cab4ea66aca1d6eaf9678cf70;
    localparam LBP_19 = 10000'h150ee443ffd3e2c99095656712a0ec771ccc1bd0308fd5da1fa817741ce88b2ab91ce39da63272d3c557e87699c41044a71e49fe9854fab9d38b95aec3fa25a530b9b3a63005e1d7cfc84ad0b1c59611552c998574b92f71b876303f7dcbf4480bc447a1b0e2ba8a3c7551e0b755590177ea0059cf49f56732c25ce3fda4fa9e2b3d034782b470103008a0583d50e3922239dddc28fa58622a6332a7bda3372de2c654c59dae3f8d7c4bc87515668ed846b211e93f1c265b411d672354b8f14268ed60ef3c578804ae58163c95b60e204c8dde62768ebd5d134c6150df2d401c3b1c079d270da3ac660c7e189b24abdea43b8a038cc6ce61a1069f328531400036c00d4d496c677fae86070e73db72770e9d09071a9adc218ba52f8572d59481c7eaa45148f18eaf522093ea34c03fc8dd750a475908cd284f9e695d0a98f0927f6644a33e73410d5c71850c08e88eb74cb8f61ceb6646b166d5204dc0d1584a8e4fc7ba6b93a2f6868d523dc46ee472f92c5b94d00a9fa2684cdd401b17f039aecf7520b645622f7079ef769278f4e62341262685acdb8021b144ed60120d0a24d344138b6c6f1ef1861f5da62405fad561220aff428eca2c7317dc25ffb76657e55fa89508aa53a146630cd59ca7c0b8733fc4a072d3f2b921eb8d5a2597fc63f58279689ee78afdcb40c1ffad6b1d50e45d6b5ac4d6df78a7f7aa93aff4855584420d4e59ae0c2f1d385a6313d020f7ea36d1d97b9bce49806461b1befed33b4bfbb7b697e7f12b2ee95295a53482274b146d9fe0760b828006db5709b47742110c28a73f79f6190fad82904257858b7ae0957371acd3f2d745c91d2df4e4e1e3dedd21fe9d6ee71cb19ad962527c3df30abc7966f5e08529ec0bfacad8b7cff0b5ccb9d719be4b2cad86e02bc26ae2608e2cdc0456853cdc402a000da9bf54af7f89dd76907235eb4d908a78d9e1aedb9f89593809e4da188af66475ef42c470bcb90fa848e7711f54fbff280671471623fd646241556655b161834b7fd1ace8169aaa87d02d39fac938317c670a45387b738421bc2f6efe7b3d9a3d705647e1a82555e6bee96878befc0745f1b11621fe995859fdd9a53446e841ba38c115b6fbdabb3c001289a92b76dd66fa140b62a110f3525abf946dad929b9c7a9e92e6a15a98b8e4368aad549dc33a498eb599e13bacf762cd861c3dfe3f460ee958a380fcd2a8296cf8add0bcf99b99ec6abd53c58d9ae076527b9863166c63a4f32ed0fa16ce744756bc30ee78a69e1a8329a9748eeaaedfcf48bd3e22fbe07e6eb5bca25d0647b4d2702711a804e8f5c63b21ee3684c8dbce8cf0427d6c7c11fdedc6c43d738bcda8c09a47d52a561d7405b738345ecdc346f0ebd95d92bc01f02747ef3cb7893137912af8aa70aec351c11b746dd00c5fa4d17137a0f306a8ed18f296e3d6d87102960d8877de34914707b02c1e7e77445e3a46a7ef4ead17d2b11e6f97a0f33d7857b7d1e249ce2ef70e406554bb4b7641d3721fd01168b0c8855471d26be74010bdf78d6235f2555243ce958785c062bdf9b243449529524f1195e918dfbf6dd7381cdd643e5c98c152e741143a57b3b697662b21a63596f19e4f35b0749ecb58d3cb87a75cc7e65e898a16809226cd63cd6521f64339eb9d2117cdfc3e4da13719a5af5adc3d90b5b45109cc954fa1ca916d7377628df4b1e6ba3ebd3f5f055356bb0628c26c2586059fd041ece238dc65ddb5ee4e10dc190d;
    localparam LBP_20 = 10000'h9229179722ea41791be0473034a30c5d20add01c4710b6361682c58ab90252d02ad3843c56b478a3fffddab9aa8a7cf9826f41b57e59ac8c6c6992941e4a84eca696fda9a23a3c5baa4fb758991afbaafb2d08acca2ac74a968b6a52c356b5d214ec18513bc6da5ab962ae3c6b4aaef4c0bd609ac5d17dc9adc54eba32711a544b6575bd797a32093904dab9c2b0a9c87a184edc47cd9004ad2dfb803f2c5fbcacf06d5f265e2afcfc8e0e91963686b4caa86262809c6d954a2cb81ae85438ce8cf4c769c3299fe29ce1b45329e140d8971a810963abb4e9d8ddd2f8bda1aa26d4609da23bd664a5caa5329e484d25b9f32f93e1c2d0db50b521271035ffce55bd4e991cca450e8496687ab3fffaa5d1c18cac30a9a56772208e4794fd60cb9b8cbafc0de241ef5ad0e521b2a17d4d5b79aba79f2ad03013bed45225fc0c4416f8c56d4a314074bd8a97bdd7d8cfdb1a9e3f4559f5f4cd0be7932b3bcc26fb4af44e289f2cd9093d74cc9f0a0d2c4d92ddf8daefba23991f65ec1df5bf5d49a98d8e919a8061820adaa2557420341081c2fb8fc7bc62fe675ca458aa84984ef61d52d793a6b80c1b33945e429624ab0ab45b6abeb2ec89f25fef999ae2fdd1576dd28a784e1441cba5c080771667091f3368e120e8ee800267c5bfaaeeafc71da9f1ca044dd858eab2e55d5444a9f755811dd5d93603d24c2eab6cd35a09f393933f936d7c9a034e6fb3e04182757f8475e7bb68bec2a9496808f9751336ab2c1f5025874be9c3f2a16a25516b887ec29fb2bcc1ce5ea87a0ad049343030c0963a37a7e00d0e0ef258321a1acf035eb586146045929558a767d183e310cc66046a592037397da78523b0c2fe262429b4fea3bef0ed35e85ada00de999d68ce691572047d4073ad3265cc6ca6c5d008cbecb768999d9b43a82f7583dfea9c37189d7a580bf75195f32df86e303e81a35e44790d39ab03736ca0bfbcc0ae2de3943e8e304e21470e08588fe62c5f04175ab93c9b178f45a21e92d6762140ddc1fc52e9a1b29a134b86bad0dd69505080e8cd641fea67fc152ae9503e04f7d44a7f50f947b9d29fd2d3ae38cc2799570c33095a224a2d7fb890d2c8eda087e5ee0fad5d9dc3689883d218b3f7e47df3ef250316e61e43934d07646f484ead184f39b1c343ae6fca5d89ce57f3b7799aa9fd38be0d1f764d6a50e204a48fbad9758b3f3f6a4295a083c2a7314235125ee6500d6085a31ebd94607ca4a4789d9db2294be69813f4773d88a3a90f911dbd22565a2ec229c01842a2e4ea4888852ba9cfcdfa71ff73005c6d3ac70a611ddf49c8b689daf0719e3a56dea536e966f2f17cb3b1858203ff4ba3f64a5faea8979962ccedfd08d7edfc765cc3e7da72683302d1e6381813215879bc47d52655bed09648f7d42e9ffa06c544cd5f0ee5fdf2f1f9a573c2afc1f805bb14e3d911252c7844f2bc45a54bb2acead44a339d11fc58cb5f2c78f674f21ed5c648f4c5ebc1bd30e4eb2fd1212ec077ccc9dbc832578ca98859679d1c979d1b6a7fecee76ba8b1e64c05bb6f49a0137c71b89ef2ee50ff980c3bf55bb2a8b96d1d6e1551bd6fd12e0d1f088d619fac80717a040b5533469372f06a0c23285c2cecaddfc5bfc8abf9e0c2808bc02fa480909b4b09db630462a6a34caf2916ef7e64376f922efe9ac883cadfd29650b887351985f83659b3aa662c81e0375037ff6a793affb43523a8db04e92815f990f13a98759682dfe850b;
    localparam LBP_21 = 10000'h93eb8a25bac2f9318f5599ad66d74515c8b2f57e31aea73cb7aa3a481296ca2f0ac1507935b0e3bed96de5772350edbcfb501f656922e02881b622f22fff2709e6b2f09197bb7a87120ea8eddba16ba2c433e89824dbfe0badccc6f9dd09d574f6addc0b4c6d575669f67fcfc024caffac7e3834d1ff28cb929b3cec151f9d65570d46d48859f006a416d246f92cea0fc3cf718f6cbca789f104cf306de1303c647c6cdadbbee2930daada3e133e84c521e34ea8bfdd85312a8baaabaa8f808bc8cefb24923c69271b6b0e14aa1d4a4fd82b793edd7489a9cb40dff28bea4bfc056cce824d6303c0a3ebdc6d067629ab0498acbc23c305ffd08ac9adb61096a2459c76b584654b90408ea92cafdc554419c93dad12ec40cded7838cf865d70ec41034e4baccc762d525985bcb7d1cf453aaa5109c2a7ad2118f56807596b53bb5d99209ec314c9a0b27104518e6391bcf9b60dd86d054232278052df8ce51fa7ddfb73c4a014f1e56e619e3a68bcea40b4c342b69021f15193bf61a3d48457e36a2cd77853bd662ec10939a819dba497e8ad801db3766250f2475257f786f49b4107ee5795b3a5063fe6224c9f842875383c35019c22abaf9d4f722bf916333c0f7e4b2d218ade37bd29af7b991dad301a86431c0617e95f174ca6c5b51f208e5bfbe5c9ccc60ff3fb70a52e2a23b153cd0633b255269d30c38929c31aa93a54ba3be58812bf2fc70bed7b10f03750cdc059b4958908ee4e2116ccc64eaf59bb3de5076e2536572f13390634d2c7368e9e1fa1067ed384269baa351584da4827732703581e4e62771e111259002dfc8cb754e3809c6a4d29434bfbfbe7213187e94cdfe425ebb66a20731b7d96ad98cb97badc5d9b49854cb245746be4408b72c16437246760022b8046806ebdf7a0e2f598974e6bd407cb1036117cb501b80bed9be5ffa871beecb2caf7a0cbb60a277342896cdb2a44bce83829bd8a4cea1fa2535df4fd124aa805e63762b3ab361a35f24a5eec17c30dde25ee31cd3d03cee5b9c5e9148dc922ce5e03100fc82922aaf92cdc4047981301f15a7ef5b1b7386ec95a46b8bb7f7c0d70bcc24738e82f02d398dc3e423c73948de01b251d234fab1bdd0f6deda49b153dc4093220e46c9a5a7693c171ff12eae444c6ef58a2fa0ad90f286c20613f558d39f9132d1e0cb3904e6c025fbfc40309ae6404b556936630ee5e7c67155b30fa96e7ad718016adbf65a8961cca7b575ae7f2ad0fdf47502feacc6edaefeec7a6d835bb22dae4ed55a2c0f456516597494d7348493dab02000b234c251de000e1ab0dcfcf1bd74918c910a1db8ae6e8a5bf4977a60d9195efd93d08837645cc748226c7c4dcab92c97e974974805cf67e889055f24460842f2667c2530e1d76040c51cfc652b0b71354565e6ffbc496fb9d61f0e74a0f73fb02b65e43f49830908acfc1f87e9f66f98e894dee5bcdd12abe6f3ab3b01d7835d825ae7327f3a5c5b034d4789128ceab3fec89e2f4c4e725359552ed23d7fd774efd6335a052b4bdc929b2fad61766799163aabd1256e8b2710e30dfd2da5eea915d434f553c20524818703675414de21810616e8613a7044955d279ad4f7e5c6ae6db669bbbe986a00d3ef85e3ffe25bb00eaa7ca32e2c072fa153c8f8490e315a765d9eb97eef11e284dc782e1d2c35940333455759e10c39943d2ff0df4d94ad88e2485a2aaf6738454a4515226aa042e8e539bb151cea226f1ff765d070a;
    localparam LBP_22 = 10000'h79f8046878f99fa7d8b970d98046c9f37f9590fdf262516bd10a7101743bc1318293b1be83674d4233d6469c757cbd5318bf70ed43d0c48789f538596d901606d6f922e61866471202e97748680cd2be5afe20d779a0a34a443a23f096bc160093bda4d9ab83c66043fd8a1780de66e9a10245fb1dbccc3975ff953b2ecd5868470f6c568b955a24b0595f7314ffaf85960defb1c1f82ee6b1a14a46f9ba493152cb6412ce92ced0ad329923f82e7ca4fb2f0a723779ed6705007a4fd2d8ba4cee56b3d522478325bf2f2c89c5bc0d23f5542d475e56f1e83a8aad43b73d18ee776023306cd410352cb757b18693269aaf46505392a5b9861ea4d885948340b6fac1daf6a9102402ac9e339992f4d56e1cc1d8eb8b3ff9e08ede238c6caab7339bd4d2ab9f44a22b429bbde4f2b9436308c5d18a526a56a5938f486173eb2b652b48374ce3a282df7fc49ce45cbbde53bf9dd393059f5a475b1f6baf2fec937c19e16426585aebc7f714a257db407e76e38d3d1ee11b1473a7a553f7be88f2729ca6083b9bdf0e408674b5b2aae9ade7c7ef5219753100a45afb7e963e076fcc3549b5d22b6c199996d5ca5760a1252e0e962c6b665958a9010b1719c11bb43af245ebbf37c2d483b1df76452603402138ad4a0cb08e9eebd437e5383bf127b50c4b40908861cf2896fb6877860062e921462aff48067d26ec9ee72e844b4a199e3c0826c3ef90bca739b21f75223ba91667f32f279209bcc780d335b35896c0897e6ad5c76fce7ce408055c68958de1b663fd0a886932bcffc30afc5d446d7b435778476773c11c041830be197bed7665bd4182097d87c9797dfdf40bfbf7cf59305e101aaed80270d031109cc2715881149c828fd5ec1b61726bc85ec020f6be658b0772bd20f1d9d10f956c8f56fb5478255097b827bc4b4d202da7d40b000512e0f9bef33e38b934701e0d2f83a2919f802dfbe77ee1f67d38c7eef8ce2d0043fd066162d0350d063477266d316c843c20ad2b20fcaf3ebfffef8e2ee006cda43f42e15feee3ac311b974756e4a6ee02944815e88725eac68078833145ee3c4d2612f1fdefbb4720684a784a94eaba38ad1b3ab03a2e84ae50e3cbaf859ee3c0696435026a550ec41f53ce3dd57f7ac7a181dd51137513f743f8cd2c6739f8cc800df4311d53787f967f26a4eac6d4ccea425cfda5cc98f2e216ef6e6d22da47667a565042684c9e6feae8883b3aac6e920258167b479419ff38ed3384a250b0660389a4092a458517df9a7eb53f651be0f98bb2dcca50d8790001d77ba032da752b55b258dde0088861ed8420e5424537414fc0775f5beba3a2bef25cad47a2269c87b0f92e0d48d67ed4e77e5eadb337ef05971fdbea1bd0842167315b5229f0f74cab80bd386663ec81233cc68a9cc2d86aa0bcb3fee43b1de33e571e125e947a62f5676e3a17ad502c9b752894de700e0a9e86cc5d89cf098861c83c4569f57fbdd1ed775d0b9c8affca5bba05cf6a6a8643b095e032b884f2e013ef11d0f719f3866b555f7e6d58321412f5b817843d10fa08963c949c5d01fe1162b96591d30c4f6696fbd22731a39ff7886fa9384d7145e1d80f27f737fc68079201a097a387a60df32f5cf63edcd5f251f9a31611ba0b803b8f197980df3275de37358f240c83a16f612f0b1d66e09959f2f8841efa180186a1415af7bcf93bf8443e277e2140837a48d7a2ecc45a1e5cce9a8e1970f63dd070ae3e45844f69db9298;
    localparam LBP_23 = 10000'h73c178953359a92a6b6b4edf49d5b21d1546f2c37f7d3ee0e2dfe480e9f26757a898487839d369e8e66a985b0596bf0b6f41d56fdbc38bc5019152adfaf4a17c735df52fba8d09eb1bd8acb5112b657c359e70001bf9fc1cd1b337143bb46c23fb036db6863f9f51a37565fb215e9063318358e70cf7e4bce657fd3fee93ad025b96dbecacb5b15ae386be97a912ad836a68ff9122d5e2792a6a6bfc2b21efd99765a5f82153cd801e26e318c2e9e24dd8eb89f03dfe53deae399c090fc85a23d7c0626e77a7aa82a0b235fefca6f46c0ef3bcd413aae5059920055b7c6c4a8b6469b357cf359da5ff1e2c2eab989c4d406a38fb3dc3356b1ef66f2125f4726a00c81e2130cc24279e50be4462becd44dc59397361a1fd270c28d3cb2af0ba25465b6cfc549191c74f56deb1d3bd85dea2f7798d0d1d2097e84093dc66ae1a53fe0d5483f433620b471cd8873d163d80c6eae718c9159c27bc665dd9e120765e440d9c717b6745cd22f1279ce5c0c873a30cda8f654f3dd70d5f093698e3188baa6b7c7933d9e2787ba42d26ba7fbcf5b8b0f53c94753f69c68e3695b29fe382ed657c19bb988a7a66b7198fef49a257b240c16c261f273273d57e43b1b30f742658c721ecfa2043a8b5e0ad2b7ae8092abdce8bd0a1e6c9f1c153d3348597d613048c9a68e42a3b8442651ebd2c8a02ccf6b09181fc4fc1067b46b3e3e252ee2d5b8179796b7226c26af0fde155bd558aa30ec16bd68e7b0bf625fff255a49971b38d8bad7e36fdc284b5e3142d6f9c5c22c8de13855b9ccbf0d6c9ede09ad25a8315332f8ed5da9cf89b928f7157a03e0790b2a235fef360f2e981b8501c916d5cb3e174e6c6f826b4440c6256097a009674bef3624280cbd9529e5fad5a6d07e0d8f1ee9e621ce2b9c4d9141e6eda80e4b79b4a18ea73268b6cb6efad5ffeae1e046f85f91b8df9bbcd8432e73d534351ee3fd8db0ebbe42c9a31e354500fde474cbb6c3e7560b340c33420fcd33ff52049597a422027a90645861a390a441871b8432d32b1aabcf4e5ffc413855c6c585867f08d0a18281117bc8030305434eacc6ada7492ab107d99f7ac9e45e3d88e85a9b6e36f69b8d1bf428cee589aa90aaf2e45ce11546c4c4100eca1a11fc4505711329ec66035ab852ffed43513f57ba479bb2480bfb1d2e83c6929de525acb490c83f59949026d86f9740f515e8344790c6ebc9634b645e3b603fe3e394ad7d29cab86beeee6846c8ec8265d79b2c30cf2c4a8a58fa2d0bbe114de882812afa86f3a98d0b1505a186c4607ab8871d2ba376b00afe89bfa42ba253e6113a63be9a8e4f4bc4d0a3e4cac27b8407fdeb4506b8ab7aac4c0faea2f047c9fb9ebc9bfcd83386340e6200d561af39a4a51c6c4f82ca078efe0590df7a9fa3c4cc52e77d0fdcc232f41604e871f489fcef42079a6ff18f6f10b911c94a20be03840c791a184c9d525b44abb7492a9c98221a725dab5026aebcb4a6b06e70cc0761c2b401c92b24da33c457129260a30041b3e1bb56459fdcdb753ea5078cf580db03051c52c61d02630f5574f7feddfde7f89e59f0a596f02d0a1231f8876c5c1fb858d42e6f65e84542643b340a2bd98f948afb334e530f3f7a5c94eb19140ec93fa5a3c227a84e6305e2120c226617bc5c4255422dca4cf7a0480238fec89ebf5e8269e0c2269f316c9589ab7860ad55d84f735e429bcae9fc1c7e410d0432b18279571c5c03420bcc0a2f6499b51c47af2;
    localparam LBP_24 = 10000'h481516a6563b997aa64e66ca2b55824e89d56a762537e76decafab4238750c120e911dc681a76f2eae1330ee8e2a90392fa6d2529ecaca04483bb199c2ea6fa98c2a91273ff5578bf264068673a278c8bdd5b319d03f3f06683720d43c459138bc6054cd5597c76d7d834ad1111fe5bfaa4b7e5949a8e1d5a2684f105a66878fab878fe209715777041f734950d7eb09a02961f09beeb91d98a2f95647e01d75b8591d222ae98e7723d11133cdb55eb0b63a5b2313daec6e005839da38149dab0b974a024f4c57e0b43cf3afcc97770c7e49e861da08f0481d97b4da45d9c9ab0aa8125357e5f30995638816ac3eb13a21e0137cc3fc81e17ca7d8a4f4c5ba341c2a9f3e1ca0b9efcd3bf2f20fac0cb9bdffed0f7bfd9919ec5c0f4126e174f276543cf8192ea5a18e944594881dbcd3e985f9e70d47df03aa975b5e77af8e554ca737647d156c468c1eaf1326b93c0897beac11ba07cb90495f34e243f4043089ddbf01e33b65ebea46d8846781fdfee25f2e7ba3bf6cc60dcd262d5e168978deaa3d5da3da51c5fa69cb3a46eaeb04905ac0148caf3fa6999d2afa6dcd72b6c82516ddc75876dfff608f8f3137467c5a7f91b0f46819a2d4429b916203fb52927466627d1fcbffdf8f305366e0431c3c61484a96cc27ff6bf1c616cbb79298d7ed41c42c9854f1e57d0a9aa76e629bd42699d76622f594394b195d61a3605b639a99fea411d4c6368620ea55756fb2ecc043c4b48029f77e8b1f2482a1d60a0eaf6ac19a51eb070ffdecd5d4ae89102049fcf81e6f164a0c92504bbb398de01a2c77f835185758f81c6c7f26e9e47f2efd30f02c75f643196d0d0fee8cbda8247d32866ec0b344996aa6ceb95a7de597e65e0e027a9bf5a3748b2abfb1a05a297cf994900305718a51749c8c867a4531bcc6a03af52a8d52b88d85fc2312f9c0695441d4afc2196c31bc7b9e892816c2388de6b129c2d57e15061626105964eb9013a18c0f686bd3e64839a3c23108041a84fa571d97af518e2705af62cf7b67859be9decb6ee2bca4717eee93c815df53cb1804380d7047a955a2905913dfd0bd86aabad5ed04272680a6cd7637a6251020b6816acbaf10e363f0b178b7bc7809d3acd240b4a99a3b7d8cb501aac551a0b2a1f5bdc5c2eb759f7a8c4c47e77f744179ad43a77dd131696fad29d58e1987318f062621d43b5633cef213ed29597a27f31b022ab594a3a37b2a47f190bc5969f7e35f412b31664286e5c2661c34ba403770cf91cd2092711b12b67d883215a396cdf884dc280ec2270ae0176bfca55a6feaa9423906c043e3921e63a7e4f4e602b2a52c85b5215e15974c82eccbc4b53a4565fc9686f1682c4dbe44fd210357729da581b0b2a30376ac3c324e4006e70eb6e2d583dea096cee4f6c3f50dd20107d5e83145ed96a80df58b42326e2fd36b3ca82364ff86f80211df9da9bf1ffcdfc10a47d42f4cf74b62bd9019819667e388f3d23218cbe74c1bfb1dca6f875e2ffd1586c7379df991eac74815d3ed6e715736f2dac141697c35793f26dbeb95a9b89260f8230e87746f83490051e419a8dd1f9dd9977309a7a9c749ae90b6eed44dfac8ed58609c765b76ec5aba05db20454b186d30fed9e4cbaa3ad65f148886c9bd4bc74cdeca62338bfd77a1290eef0b6f4ff09328c506d998b34843c59ad21a51d217a8d12e801283239885995694329b4c5c4af11e8209c71cc2b74e3eae48ff272ffa1acb48f49d23a2ddf2;
    localparam LBP_25 = 10000'h6f49de8d73e67dacf60705802f0c80d3716d87723cef1689e101ffd4f88dbbae1f7c8d91c504d2f95d1ba857f2a6bdf8d4da4a7b5521f321de9edc0177076745c600c01f6ea97dc251ea91b98b2ecc88c460d99878e1af729af295d92443eb4feb3131f2399512bf978dc36c4f94ec5ab16e622ed0daab10b4b2da5b2cbe87283983fc3e19b6d265054b6e61b45133befd0ebd0358fce5063924f954712179334f9194a7bd1b4977a90704d6ead71ee59eef8a104da4351514675bbb0a2dfc6abfa525333430bb754242291a8e5f53770830bec5ac29fde2a1e44b5f8e2cd573cfb1a281b0ade89f85d5ea1035bc5eacf7bf596a8e04bdc4d418826e7b9b052d2a751ea4c309d67b200e2942d27b0630bb283c68a854cfbe3c13c18c91ea6d7b3cc30b7c82fd2e1f67dc9bd40155474f3db0c555159c032d3c1e39e5ee9cc1f34007d7c0faf3ac4f1ab3b0b3bbe9cb61ec16c6b5c9a0267e400052a4aee25dd2c8ada74b33f8aaa65446e05ef800cf33e780f2e520c52a3604679027765731037b2a1f8f469b86cedb33046ac54d79cee71a24656cb47dc6e14da414b41f694b65ecdfb99c33bbe1800f1079ac56059339f4a565f42e675eab11bb1a48e16f99c92562cd66d16d280e72ee173cee564b7684a7d3520a9c84408cb5e5142cd715dfc097901e15ca7d130ea8dd94952e7362f6aa3e182d914aaeba8599cd72ba86b3756931c8c5ac872bcd947a9f9869f440213db49a0b3d732e8fffbca4d0303a054eff049269c090f79157d11abd03d3aaf9ad4da08cc9fd35d1b441de03b3622a4803f01ecfe131a7dc98f7eacc9fa8e6e6e7d0ecaaaeebb99e73bda9e948aab74e3a14bd532daa9ffae2091dcf2effe158955697a29124865a8f3d400ea6bbd9dc5cd4868b7fa31ffab1687d538c0bccffff087242cd20228fcfc375eb03a05bcb59dc8e8e523f68eb073b6dd316fce48f01f60a11298eb5144771cf4460e0dd73108fdc0170d5930927644e2b454219f2436bde4c5a4667283ddb86df68ea035aae18af75e8ce63c62857db958dd5342c0ca2eaae0854442f80abea7359e6ccbc7c22aec0d2c21b1f2c16c357c193886f4745fc52ad83c613c49ed47ddaaf7a917e60409e666cfa77be83fe9f830a83db70d29fc2990f38db22f1afc9c4490a608557f00a04f857cc945c267b7b9dbbec8bd02fecb3368a4aa7c84cf0691102548175c60875c68a35ac22f8489eeed7b7703cd4d53285672b05c1556d2c0cc7756cedc65f315e84fa11f01f165fbec9041676c48791b6fc8144f672a8b55556f9fe2823a7c9fa23a68464a55277805a116df83ab5ecba49b1014766a4e3b0ee3e5627c455bf63f807dfc08e345f5eb3226c7057e98b6c07a651fa5133de8ae429ed4e9c32f927e91e8101d4a0c2af74baaeb86dbd5f23a3409ac86f1dc1738dd034140fa4eb17143d19c12de5d0ae8cbc47b23260538bc803eb5a5c5d37c11a40d74d9f185de4c98ee4b293ed1da2e58657d7fa66e00105e9f93135130cbaea224d7d31127306c24dd5881e4067141dfbe432122821cccb6b7a0ac6b9244bda3fedbc12d7c760793271e176e4eb309176293d189df8e7b39a149fdbeb7dc750b2c91901a0bb7807819f792b200c9a193fd8d284c8971be3a2cb14b490994ea2aba16b89ced999a99df8a19403697c24eb2330683ae1f02c6d1ecfbb7abbd852b85210736dfb72c10112ba1587a47910db2bbc28286c4d1291d6dea87dc97d9a70;
    localparam LBP_26 = 10000'h8c8483c8cb931aaf72bc9dc8beb9adf7ed062aa64dafda32f6b6644b56ef4c100fc1a85d4b0db986649069f08ec0dc1d5ae0e17d2c1b1bf5341bdd6982f880d9efa0e11342f684f5955bc9ccc570579448b8131c8caf77c5bcca2460d0a1a5d1d55ed20bc547ab8ed755a282fed22755cd1d8ea93baf6cbc34df4b94a8617e58ebdeb4dcf1ecf754c9b291ae64f760d013a84306d086bfaa308dea8b762ece03072a1bfcf024bcdf9b781cef25c1504ec054643408438a87013d19576c82b95edcea6fad4990411aeded264f1e15c5365b98135887aa3a57667abab4d5b2fda23bc13df62879aa2412191bc5d50b5ce06c8164e715e63c51381912411a3af6d1db4dffcdc97950edb8ffdd6036c83253074ab840f3c317f816e691f4e4fd154c1bfbecf8a70865fbd6256006aa9fe909aa118efd09ca741fd9c678965b3b9780561777559e1308d0f1af35cec0e3febdc69192d32584e71cc55cc8f72e7ae069b7b6e29698b73b17014ae09368b01617a096056c62d093dc766d9229127066949009e9a9a0b7a806f62d65350f7e14dc5f28968508abf37d13ac5ac412641708648a4a0d17dbe03ff98de0ab9ea299bb3db30639bf632defa1b0f696a2788ebdb870be2a3a23529264758c986bb5c15cd8aa367ce7a841b4fd1cc589a951defa2b5e711b7d0c65b072a8c44a37bb207b5aa2fd75b708d5fa502557f8662689a61aea30ce2244e546446d6b8a9daa52527b3c3a8a340a9625b7f659ef9e8b8fac24ea45f867997a514092d6d29e49497f10b3b85ac28fe6aa9da192cda7561ebb57ed62ac9b44a3be503745aa9f550eed128f077ef9f42f64a8fa7f6b7b1114ed0c61d19425dcbb9e483742768533065f571634ecdd446d64dff94beb90484463bcb0956a2e9b04877b79a9a1f68dd9a5d878adba703294cac0a885823bd2386febc2dc34c64253f41163083ad74cab9cd675f20ef46d91cb9bae40fb1e769b6ce6e9f2443af816078b8f0bfe846283657a8594e22fcfdbe52e3fa4488993159be3325dffaf6c260972c650d8bdb6fa4b92d8c76f8602ec7c7a355e6a309e165ac6a9311821205d73c395605f308e7d5d6fcb6cf7970bb79e6a0ed8644baf42520d1cb38b16e309dcd1a78f3b3190b9909e44b6e296235ab7d39611b01d0824339a6e52bdd7eb9e48a3322bb260c36326e06891f8ac57f0745b6e8f4a23075b1b5ed215a9f5fe0b64c897c15d8f136fc70daebe8a96f12d8207973e1ff6827f7f9d317493f8e2315cec6979350a3855ac77380cd42038b0322e023caacd6ca9fd8d106d26967e4e10422a7e27492593ccb08194495593970fcde672c7fe5bcd384516e5da52f3c41f05609c68e6765c8dc32e8d9d4e5fbb8bcf162594c912e3325e90484b195645e973cc14461dfba7192970352cda9e5c5ea7cb524668ccaafa0b68b1913b8e88aae83d5e322149b2863eddbe076034734371ce6d9d754d3662a25a4e3d18762560e09a1a69ab471a8d69aafab0123eb3ca12e890b42bfd963566a6121b2e2f4c0083ab11837e340084a56ed353123d9833b8281fdee3c85f2723f54d946d5fb5f7b3c5da7d30562a492bc8daae6d78ff63965cdb8f4c8b05812e7f6eb1b91686ae59bf796c3bb60f25a54ca65b0ae1b84f23648c0a8cfe0dce0b05d1b5503ee20b20b4812211df1442dbee59074036997f1047c29081315c200b0f4d170f43ff7d36d9754a3abf1f45f66b3f90b33cfb8a24879a9cf66b42b39792;
    localparam LBP_27 = 10000'h1b4d4449409de82c2984b7f4eed91433b2e5335b017b5ac103da93b8b79392d3ebd72e89a95dbcbe5a1902e00622c1e41e69db9d1ecb0b017095b10a462d2b6fe81f365e690f64f30c43cd9beaf13cd001d474bb9669d9ebe4509f24aa20cb0202b682fc31b9a7981350c9e20617f0e39f90ff26c6f8c723e17a4254395e52a73367c8593bea69e4df2b871e103b44d4d74fb965b3b1ebfee8d2238346b15d7baae1610ba6e67c424ba7686191acc3993cf7637ce4de50bea71b90a1645c6273ff45785b3932b4086c9784b5ad55c80ccf213bdc201b777327ffbf8e6311f18178abb478ea82733700638ff94322c4e6e232b652d493ad9a988eb1346d8fef8f7ccd4429cf34f7690678ace6bcdbb92605288ee9addbd3afa83f22f48d3193de62e69897813b73b230611d20d27c4af3482fb26b7f4c40b0d574f6de837476088f7536141d7bf52a217a735a48b182292b1e14530da97800c48871ce094927b64dcc88e13ebb6d17f2559e2cdd29912858663eaadb9673b5d7d1bd6729c92a31795b072ac0fd0a236878e9abec1a07f801c9cc0eff3c1a6d966963b4c22a01a1f1e53d7f96c89d73bd9d9cd4b42d8eca4ee043bb9f076f21408e25646e0d628ec7c88623f5d0c3a88613ad081923ca0187ebdc6947369fe3be804af077f87fffbbb2de4946f268ec6e07cd5067a5a9ff7e9665ba2967bbe0012d36e8903925e7cab0765daa15bd0568851440ba1a010e6000775f9cc7bfef819ba8059ebc2029eeed11a2996baab98059ec734d75ffe4cd6f1f4a687a89d231d803acd54622da6af400f79c9fd05f565ddd2218c4d458ce1b73f6ebd1a1143a82d8c21465ac07708a50d6ed7ed2eea9f2842577bcf83a8617f4a3edbd0c58a27665666d3efd905dd0c36a61cc7440d44681e487a67b44b91fd46c8d267ad7a54a8bce9d4743420cf6d602b3aabde6a515dbd431f7e75005e88627cde45f0ea356b47f70361c67b78cc4e1d841cdb8d0cb0b85ef79184f9f55d7bd537edf95be22c75a0223b1291170f821e4d4c83f052b47b0cc00abf9a1bea2c4ea957f0187794a12be953639f735028f24b23534a4706f461651dfb09f304f6dd0b4f0f8f1c810a5fe0ec5cc877855f567a082cfde2bc2c9567bdc278c2fbfd96fe6521f67f2386b61647cf2fed4385e8c0661d94c06ba11ba1e49b52177f2f05395b800326aca4290d0a71eb98d49fedfcbeea8da0c378dc40088b9a7afde05a4630978eea8d58c34518b9b9c43f17de66e25e1652b3a186d7c03c54766a24f280102813a0ce399781dc66db31b9c59d1a2a892786c17ba9155230fb6347f0617b74bedff8c1e8b027afd813ec524c550f0e3be38d9291ffabb035e9459cc92f3f571f4d4344cc42c5edecd7397ec29386c4c14f7ebd2effede8a1c1452f2e2f7324cb0c76b810df3d374dfe0ee5e539cfccae9e671f76afebef2824f137afd946b0901b2b865862046bb01960302742dccfefdd969325445edb49e63259bb80f02be94399e72ac2b8de9e985a36b98ef2cdc6c4af2c5f90afd50e3054e34ec43215205ce0b68f2ac706a90b822ab3e9a19f3c6abd09cad8100a4610c30aa9c3f8e2eda753de8b8ad71409f795983a3ef77fe516a954aefb2e58e417b2691411f016a8bd0f11d490583dca622b3df9324b8fa05aae4e9125d1f3a88ea6b488f27dd89e534901631aefa53e1fc4583dce1d6cdcb099e8c2892d4491aa329115b7369189029640064639260099212;
    localparam LBP_28 = 10000'h1f455d7c55c9741fd427f1ffa7d239409ed6281ef306e21ea5107a735110699c03af3ce765e07c3f419e8d6b52a42c25bbc5f5385346c25d1bba4693f0e70197b1d2a5ef474b029e975daa9bf43f5e4302bb01d020d086b134e4c08a2983fa0ca0984529b800f89c5f6d06321abf27a985b851dc1a380326f4a36cbed5a49969eb66532aa6046b0291dfcdf4413c2c43ac12c4ccd1bf725ba34817e862de93490472e98f30d18e92fdeb89858d3d816a0be7eb926fcc4f0a9fa06b5efc2fab263445ae28842af2e2cefda5c470c763684a1d2b93a5060cc476dc1ae44bfb692115c6e4e79a7eb8e364dad8b13ff4d3919a302fd7c9302a6d79f98fd6a92b0a3abfb0994f5853a0ce8e417b4f31edda75a857778cf3474ec72e3156c0641a695d7cac04f425b49573eca50a3e583b052d43f2652c2cccfca8d820bcf26b1fb23f00bc81bb8489283045156e2d2a33c05236f65ff7267cae70cba89589441be712aa3992c930e3bee01c978354fd388a870ed7c13c62f16b4531ce0885ce7646e645b69bdb503c81ef18b8d695a87d8462d577af706340f56d85475c2ff2c8910be24d126052d5832f30c225413e6d5f57be2a805c21cf0642087409f2cdd6331e175f0682c3c28190bc523214a13450e87454447e7c27090048ab85e2073f135107bbe8027e875c0d5686be113393a9c4aef9f6e475467dd911e865ea248777837125f9dc772579e2c96492821d03f88409fb8d704ba8b3725396f8eedd73c75c7a209a63c43d68bf268bcbd87ef23185273d7760e0532594f5a7821f679acf59eb1c4c2c4790fb241cf141bbe2071b00a1bbe0cd3d82632e5a2379058c23e3bf8f2fb7ea962cb9f01f7205a5938348ab37919d3cc15feea202b2005bbe1e144b4078f57d7358c18c567417de7a161a48ab3a486afb4dde8ea2d1b06203b58492f9e72dfe259a71dd537e6ac55dbd815c02d90a649cec1680a8ce07d0350d900e1f6848db8bd44f729563cca57103ef24c60f1b88e2bdb878abf7b07d01bf73cf4abf1b0ba7855fb724ec2d29ed1751735b2bcbbfda02d0debe6a5778c31a4f3d90d0c2d16c85744653f4b064cb8c1dd74e071d11e99abd9a46c10f651fbe6637ca0f4766968917edb20e51e70dd9fe64e76bf5efb04f8d93352a286602d64161e4dc9c7a28702b78975ee91e1db5294602b3ccb1382f748df41a82b70c0ca819241588b322d02de26aae673627d53e9d1a7e659479590a04fc5cf5f8ee1b16f20d45d9fd95a6d5ccc3d9f6ef6c6ac7d6cd8599905e5352815e28d736aea77c6c7b240b18a8289506767ae43c0772f7ce8b0e7f9d93f54dd60a4ace34eff4ca1dbbfa247beb9a941678f17aab33b801cc97769319b4ceb6a0f5671e5fbdcad541414dcc0dc2ed5c1eb5e322e6173dbde7a82586b6638d61ba13032818f8843434de7d0b2f148a982d887c8e9ee32ddcdf118d81a66fc64c8fa8bd5cc82aa5155b9deb18a620ea6bfb7f9b0173245f53ebf83f2588fb94b9526d4cb4315bc0e83728ddfdb57a1b75191df89eb7cb51b543f432e317e9007e8f0a8bd3ccfe7f5b3b71837c592abb26a268c081464f160dbb1be49f14a21cc37205a82a683e01f45a9a86cd21b343ca1600c80e9ac7bff72379ba2c2bf14e4635289fac0cfbba27e85d5188d83aaeb8af605596ae7f756b5912657a6b955aa1eac468b006351af4dfd32de41dfacfa95def447a175c7bac8f8898fa7b8f6a495fb23a762aef178ac60b2a;
    localparam LBP_29 = 10000'h9aa90ce6c8bce87207bd3db30769937b7006831ed9c6bfeb33055960fcfd5be72a7633057a8d1f9b879787881239525fa7663f3df631eee5626a2ffdd44f7bea7b4771504b37578afa5fdef4585a57c24367add80b2e8e0fbdba20901bc81e78dd906cc83e4991efe5367ad0eef824df80deb9f4b13314ae5822c06fdb7ba2afb20ba9199ba1d2f86a24228b66c4fc4fb94e5a25b279959fd21b447449dcd342f507e3fd1cdd7c02305b725a20fa10c60733612d31550a0745e116a24d9d2c9e676f6b31f9c4e70be98da61e3663cefbc85e1f42fb8960f31644a3e86c53abaf21b4e04d94ea3216522fdf597ab03de8241240c419fb2eef106ea8e741a1a382326f0b7526e7a0af7c2f374d7f96f92ccc0c6953c97547ff3e6bd078b68f719fb01fa8e9d46de33b87382efd11da23c6c20c5305d54b4fba8b046ac8fdb3f98e876726989ccc571630d04fc52bb86f502183559acff5a597613fc071cbdf1cc73194a94daf86c422792f258cf984efb584cc8e637ee3e86327520d93f7753ea1d08edee0eb660266ffd33476daa0b6eff2048a8e1f92fd9bc64b7808028ccda8666692c579693bde5c6cf1cc2502d9be753212df688a5dbfa1c7fc2ddc9f058f6c058a9f2597f29e4fe13551429461c11eeb18562100f6b4479c1e5b042dbe6ab597d54430d742aa6528947955c9af7015f03d45a354d20333861f88db7471dc183f7fecd5053d841ec55eb675683581969f0f07da0dcb784336901365071823bf93cd928d5c8f5a03ffd976bfa5ee79c0e1fa30b538f7587f9c61356f9ec61860bbc22089afda17b308743555e182603600f8256ee89288dae5078d113a1c6abad4b26b3ae6d2764a8ff96dc930d8b8e032637b4101bbe1672d40af3c50456f5c466a471de0e9350825dce6b98179f6134141fe6ace4c69636459a1076294226c153ece4da0a13a8bf99bdb69ce5d81b7f8d09d88e3f3e133c2483441c31934a7e5f8634f6390a906a122cec2670431644a92be36a018a1c2be5c8d9b847173424755c96356080cc832be55de891d3a04f16dbb65c951e0b53f5e9ec302e3c772e6831258f229bc32495bbb9a106fd56e9ffa428c5299887c7e6b49ef6177931c9024d1da327fb3ff0624d96483ce443da636031567d7b75080561aad4322d7b34a2e191497df386d9925e50ef9d67c61d51035a61ee0280e6959b468fb00c2a789567f01c0f5d2fb87fc2d93f39c12829d5485bbd64b9ae80e91960be3caf43ecb2ccfa5eda1f03d08c8ef59ad03bd33cfc320fc75b8e0d5f44694cbb43e7f8ac23ee97f8874304dcfd689cd0585e1f748536702a9f6586cdcf04533de7f242acc108ce85839e4825489951fb6a7e2b6962119f6ead62ce8822833ca2512575614f9354a194f65362bdca797783b8a10bddea3f4da0354a3fd05b5f7936cd00ccd9060c4ad857540ff5b11d8077b1a73eb589d7b7c3ddc4893a1770a0de08dacb8daa4876f3b5b382403d0523cc146c5fa61e422651d291f1d9fc0e095253f8a0a7ed932d5976356be4dbefbc40de7934c6f802a03b8e01b11896db9848299a0aec4fa484e33579ff56afaabb0d65490e44738883044febd98fea1412162d087693ad2e8def06d1a7775d68b17b3f7d1714c95295ab663538fc281060c7f150316af923019432acad3a32d8f9448a98a28d21642e5a29aa636fcc87710d17a703823ec5594c861339e4b16e84e30bfb7aa662237c21fc7f24f13f4b932f7951610;
    localparam LBP_30 = 10000'h9f56e7e8c64124c87907f5f287752cbf0f285d3107710af6c9acb434521123156e0e7243928b4bb7adca6effd325cc0907c24239cb6777a58f4f3d5f1ac1f144129136aeea82e41bf77fad66b7b53ec6b201764c2e540f496e65674e8a658f4838f8ef89425a2b832be1e1bb5b1fcbce08b1fd2c2b0f57be96eb42b9b14fe7e8e9384b9067cda785e54a370d39ea0cb159984bec37d8fb7c169d85bebde79b4e0e63429eaa0c3c4ff8f124968f4ff5ba9928cb337db3b800ae05d223c82c4a0d1e5b634cb02519cb0ee66c663c08a5e6c81569571b446d450bc94945164a6970986a708f812da170d1d6d150d64e8ef15570393bc292fabb0e6dbe7cbb92a687fbd42a60fa7b86bfb72c84fe4ba3e88c361fca1f2b17e6237b1ac28369b6edce43ca14c162bf7d4f287e9dcc41700a87763e3e27bcde8b2f4ec3019d0a8684d27bd3ebca22c44d1f48c4c96eb531ff2fe3812fcaf9510f36b32ff740dbe5827d3af86e1ac3808c2cd6c1bce7af6f59c240a52cf78f7cda9c7e4efa3323b4ce40a1f9da8f73d3b1c750ae22bf46a6175e4c7c658949e9abb86ea79890375be61b343f4630ec756ae213e1bad053ad8422db869ac929afb363b7976a15a10fa6b9d94c287e6b34946d6dbfcc036b4b861fdef641a89eb4e6bd990afde4a4554c9384dff8dde54ea9f92673f6c13c0a59d60b8f7c24f070d785d560a52375ae9aae2bd32b78deeeb23ba78cb82c962fd90da32e3497c2063aabab0c090e2bd43a24511b061061f4b8053c487f9dad0b63acfe7c0181280edc1fa8908a12e0e249bbdf7aa6b156f0b90f6ef4eb6a5e977d640b04070db0843d8bc9dd97af8bf68adcaa2176c1dcb6e9b2fa8c050a2028919cf6013c2a6b1287f10a3a8e9c0f049945f88360b930965b3475aa907add92a0b765bb3085d3b0bfebb27c3b839f9f17520c4c6af1b2e55fe40395e615420d4e2a279c01f1a0732bb952e898e648764c3e3150ae0495401aa977a6354adddea072b83ee67683fe88a1bcdf8eea10d8b30797e87f3fd1c0de6deb77595788e60da64f195ace36068650031a7ff10b65d87dcd48b6d260ddb2a1eaff065f130fd11bee8d4f9a8c0f32d6ae21008e8926fe31106fc7fd9790ded1ef85a329af872595d38ac2fc196f2880faa319400210cb4af352027ac8e0bc023bb8bd5ae13d0875e7c6ed59a89900886bf0bca74158987cb16f6db85b3cec9a338e8d3790c4e0b1496352bd6849ccca85f2177b6dc082dccf42dee8db5cfa97df5a5398371e864b52529f71f07ea042283adb6088d0d10bf958467d6c9a626cdb90264e2c3acc70216a1ef910a0fc1cb42e006c9ab3b94150077aa51a2fd994768f5f0c0e31246d74fa7a377588e1c42927c206009f6950f42415695d82cd2cc88f879aaa7e19b693506e2e70b508c2a72d71172c458d6683e1d9f21b9cba3ebe7ea9b76ca86f092f4c5f59d91515f0e6711f5e55befdc1a14250d9c32666d03374e2bc034d56065b226fe6cbaea6c749c060af7b71bb9086fed29164618226a91bba8d2f493e6cf5759c10f083220bf84d61fdf1b66af5ed564bbb3b9d4c98d7d4cd2e8c831a1d53a91eba842653dcbb30a420495df1d24781043bc68758aa7f52f26adcf054d1bff1326a77db002ec4904d3054d050004ec8c91eb0b1fc9c5b0693cfa92d5221ef7944928c4b74001aed2c93394be55b679863828b6a77ea72eac9381dca7d6e454261156853f71bf52a2d71da89ab563103;
    localparam LBP_31 = 10000'h962fa62746f4a643dd0cbd7ccd1428bfc8211e01381761373edee0b0292a4d4cfbb0f2240b5eb53e22853d70432b46f799efb43b3d18082c4792a0f26818990989690ebcfcdad243e374e93ef92fced70fd01f831013380d26f1d75cdc9d246bcd4d9208dfbe1e6ffbc24d1f84ac5929167a49b18406a93baf48df957834af6485d4ea8eefc457703144514ee8b31cdb500aba26ed609b408e1d0a4560d6bfc03fad437994f05a4f41593e284b0eaa66007a091500bb9415c3727fcd80ab0b25949593daad3ff7dbccb1dd4a401e7c9fd570317352595572f3be4a14b0ff592e3a570cd6c6d41cfba32df24378a1b26e7d9c0664b1aa0071f61976e8c4b15fb56a78b56552263acd1bf2a57c45a08a2a489795ae2075bdb46f9ab295e530f1fd5b7f9fd6bc414927fe8ffaa3c1cbf6cd95fb6daa07a05b4bdf584329258a766ba0fb6b1ba6c101aa0f968944964f5b0f06a43272a6fdfe006f4e947bd3a42fc725fc1221e86cbb9ef65e14ac48cec7a1136c08f13a2dce755e60d90b5a457dc7a43a112b6d94801b888f5b852e533e841f221df0fbb788602abb02b65a214ca57ff6d123e8fa0d6f429fcef406aeb77dd1895513a30f1a2ae125f75a23aa4d0296fe30a6559bec4d588be7429e0babfbc13dcbfd0eef2f4daa76ab0562871d6a90589c88d08a66017ef6c36176b2e8140e5faac432956e52b9f7fcd2ca06c82d2e4ee445ea8f4dd3cfc5fde43bc30ee6750543ca456daeb43b1735ec5f6c246054ae4789ff81d835063138895a3b6813c66fae57347364b9405571d6b716c74e6b8caaa1c272b088d9c08cd9b5cab4164434c1eccedc667078f15e767938471e903964fb680f03246005add77bb7ae19ea2f5c4fb81005a1f892abb7aa251b8de59efa72e766c12874beea522e86f9d4933e7d74104813a6930632072bc6cf12967336e834e2f8ccd5a724afae9fa1971a4d3c1c234771e8dd996a40052295576ec8a7bb3e72f7a512d016eee655865f7e11881d24dbaf445e731146939676274221291d024809dc1a09fb92c60960483e7cc5ce28405941a9eb8b2e6de2da8ae7a63dcbdac3268077c2b9dad2cc114d9b37822b7a0f1844bddb69877fd9d2212e72279ed53e90d087d25f2e6dae7b968a80e332632b949f696939358dba9af3e9c23314cd4f2cd1bfd5fa00cc083536d24dd548e7a59b4906ce7dd2fdc822a916ee3a14e4a5638544b14a84684d778392a7a4a295889d375a039e93994707376bf701b098673f0b90a14112bcd3e8ef71cdceba9b8f2d174629df39835a8b477dc9e2f745cb0472ca44ab38ec718a2463287175c7360b5abe8073f69f0980ecf99a649dd41ffe41441859547e58b2408568cc6262b1c5b430bbace5296cf6a0ca61ddf118f53db205a6539fa87934f9773445f62b335f15d411cc36ec98bebd4c11f627ed7cc9083960f82688c8078e6a1bd58723436005a447b0d3a0f231b03fcfc18c8c5bad2b96bd9ec3d4cf139dbe3b4fe0caca2d5197fb5ed59c6d4d2ff0f9a65959588603d3ad27e03bd84940d76d59d0c5e1900b1b4fcb716a8a4cd5bd30283cd31753d374dee6d3665f5bf4d663ef23d80e3f2a216cef17c5015f3939544cb7a44b601d3582e358bf9ae3d8bee3fa9079218a8efb359f191307af48f9e88d26aa257cb6033582618abca3fcdffbfcfb13ee17945bf0d698ee1942e196a76eef70b9d53e707d8b479232000f974c87020822b9b9865c27206c29087298a4;
    localparam LBP_32 = 10000'h903058589ae204b292b8144f385a131f4eb66980a6853ec42085f06cedeba928c12608662f575990eb8345a80fbfedbc59da9522536a10f2880addb6d2f4321d9cf2166e325b1e1d80cc107198f45f20ee0bec76f8bb7fbd06985e86aeaaa724911adbfe0612b39a975a17494ed3847e7928322e570c465fde6f58955c1e27f61db6a0de94b0965fbb875d453aa90c8bbccc543d6ca854008f4cffacadf2184616e10f060fd9aaa9af6d108f2fd7569d843ca80bb909b4a8671b4a8ac415020eba79ebd13819c597dae693be7a475bc2232a3e75496a5d508e6c374cb9d681b40b6dba0123468faa0a4d52427800efe81425fa04989cbb7d524107b9c7c64fce8dba3ede8ed2105aa0f868a63247bff563614025502036a7e6f1711730bc378a3593256d0feb9905e50af1bb82e42505f45121ac5000b29482e50b21527e26adbdc4b85565e2eee5a10a4bb752f3a1501243199fe14b2550278e8ca976b7a6d5effdabd252f257eff7f2ca277c17acd868990ddbba623195ebe16cd0761db26c58c4cac411b740082fc0cad98d7a59dad9ffd76a58101a8e2dca775170e73bed6869b41b98b9903d0f30c76e1d02ec58fca1deda61e8a160e82bb7e006b7f248088c7f954f331ec5321e290a3830ae2ea64e03c110f81e154ac9de3e13e6f3f1bfb2efa4cc0a28b6c719f6375af91e165d6f644475fb922cbd3d0b2315e17e9b822bc2b037491d7ac337f1b604e910be2a7fcdb66170c3e989c09ccf952c75e8716b9caa7572b10d314920564a3443310f02765a2a6427c3f354d9b8d46a49ae69ab38a053a8c5b7056711e2b914406f470cf9f903b8bf326c9337f154327c7bcf711c57f39191160390f3ae4bd63df33703997c2f38b5a1cab944e6c095ea877ba5f691d2d5fbe98651060ea8a5c6bc2a73ed36b08e56279caaf4aeb9d886d3b054aa788d189411f9bc40f9656b408fff64bf9b0a8b8aa4ca16bdc558498832a2db13e1fdf712b9b9237642ce2fb8d7a9404aa533d85044dce0cb0c153db55b044f624da51559730fdd55af9e3b0bab5786426ff03a1b945d4932538571e5e86d0aba894651bc355d6a4729213d0f9fcffd95df2056fe6aa3c60262a2faefde14c45a0adc7f4b405e88f98b305a1c3ec1dfd5f4d92d67fc291b3c1e15716f3b254a2671da307484f8f1f7a23a80ceeca8a2da85f1c7d468e4672947151151fa8ceb07aea873b66fd6b4d1582f49e437c4ca56c34badb0d9b56dda870b975ce5ebd6ae13b1288153ee581c5df18ecc9781be271b32a6405a4a17723acd2d725fc553a9eb65703435fa7bf0f6ed8db78d6e223d09cea2cb7830c7df253f4e8119011fb81bb5231243cf558faf4b6810eb138eb700e130b17d955a7abab7764ba0e6431d432097dbadff31d448014d6607104b573507168dd4c0fc932781415e8c41df6d28ba804b714a034b82fc720c5d161b0fb5c869666965919c16d5d3a2b82d8b4215137c14de7f9f3e981d3a4c3f73ad085b0faaabf24dfab0dc42a0ea718cebfee92626e21085d5beefeb4a8b38c3a33df2fd6a46d683069799d8734afafaeeddc086920b0b338a47b6ee28051c79c0142d85fcdfa0f661a7ce1bc6a7209be5fe02741e4d8e487b11ec6fe2eaacfa634dbc9c85e656e4ea46dc5dca0c1178a1d67a040b726bd7d5bebd11fac5d73def2cf232551e343c5a80f46bd7ded9bf4a64ac3e21166e8f9ed788bec9fe6c99593f64fb2209c9126ed425efb29c72fd84;
    localparam LBP_33 = 10000'h604bb605f4e3d5e2aa46f63187354f02adce9093c78191f2b14dd6903e57ffe8d747a4fe18a16531047e86f11ba009c082e9c77be9baa26c53c7a12d0c155cc94b972c97d84487787211b3cae412f97ca99a877162bf74195a05ae72afb1d1bc57444f7831027a111ae36b631102a04cdc5940bc3dabf0c73fd2c6da0324eac7c141943199db159f291da3ee2128e892b2048e5f640aee0492c1582342f99835c28d20e76d85281c18b71adc76ca742a3130dd7717416c7450c63c0102bb179f4722fcf8d5fb0ec9656416169fc9db3dbd9226e4c3655b097bfd6904472d8477195315f2d3e4dd5783be325ffbe0b72e23f8541acf015f777048777e887852a6a54b4a62ce3325cd0f7eb1ceade676ff47a02e27fc9f74d64210e934b4d5dccb2d36b776f2c71efa14912d4cb1b9a05294689eedc87d9de5f722c6ac95f1cce75f5460e4bf1c4d494b81b42a77453aa4cf311950784c0110dd1361fac4f680cc3085eea658a1443edceea81d33d7cbe0114e9f65d8956855c7f00b85e1f0578f9ca2fa86e6d12f3604070dd47c07b35ca8fc3b8f7781430ea79482c0506cf30d0145798007081206d1c173fac89ca5acb5015e4cf38524fd44238641ac5e47218046649c89b76639201228f92e24413b10c38d1de2aa23b3f75fff9705af3f625c0465cf16f109743f48183eabff62dd9570492cb8e5279849e2d4d58cd985389ce5b4ead44684a78449a2d6b4145aac9b20b589a116a7bc6590713bd8d138256e7d16efe6eb5f6a0b60fa8230579b230ffd48a9699f603fabd6ab96df23a40357f0f77b528f12fa633a06c32bbb6d3a35338cbc947dc5449b53c9da22d34004cb35c4c0aa4aea081af1a8f7e129f3c651b49d17cba0791f2a964c957e86ff00b3ad85bf5f475b83f54bca32d5376d2d6920fa148470518563ed129d3d3cd61c9c57015236f08be385bf9abe2b6985502fbdeb13b9d26b42c06a17f7bbbf94cc57ccc9a6196e8be9b5cdd4085fbee2fb7bf5f7b332eacca3c5b488fe86e715eee4a5ca1d40e01445675e0dd4b1bbba07e9555a81668f6f45541cd9ffeb0537bbf4db9761c69902f03a3fccb7ffcac44b999b646a814bd0d0dd3a2be0b3d6894152c65bd3dc60d2b02a8e9fb771d15682c0336769f144bff34baedbf7f0f856cb56ea3c8ec8c0800b9835ed0a10b7dbc33fbbb3c3e607735e7cd544200949d889c2149462fabb3fc8d280c2339ccd433e8b6a7df0c94a2b0944295301b01b3918dfef38fc321cd16f7054872e1f2f9d20271e272ab56248ff67813df8f84de15fadbb4065c462ff27cb7f47d4bc97481f5b2623a1e7cf405ae2c7195560ede97e627477f6e09756a1ddd8fa03af57dda12c50a831b5f334f30aa45a90b1d38d8e238609363d36267a690c71bc6f8915afb0984278679f6a7010dea23ef700770d551e372cb866a8ceeb1e7b6ab6e797a6d895febc089e24eb473232175cd718459e1d8c93cf33db35109b0ce5482b19542695aa9f0b5ba7f770533b0ca3e10d62499bfc5776bd11c4224b883622111594f823f10d813269c7b7f45fb6ea4df6cdf157b48de5414b8bee05061bb87a1afd79c512818ebd6880661fc4ff7a6b55e7b4b94cd297ec749b30be7aeb88b00121a3c0d6aec068013ae5718d53fe3de51b2fd3cf0ca05eb76a5e12d88dd0b3ea9a55910134071d149f51d066b64490d65828737ade22ebd944ef6980ba9e46eb06f45be994f5b7047502291d8e10d5ebbd08ec;
    localparam LBP_34 = 10000'h14f7c82ba95b502531700770662270fe4f93e9a715e351ecfe492894ab42a778feea152bf73fe070d075cc4b2b1b037a04ea8fcb0b5d8e1349ce7f780e0ae1242f7c576393933c1f52715a3c96aa0514c2346b3b52ba26028a3fb232b1d4e4434667d2f62c3dd648f9b438a3f2c4539485eb9d2820c49ceb0c5d1ff96d31331d36be55ee5a5321e3363bbb0d0cc1e1d295b9c7d57c3e1d723d50511af6ec63a48cb164412697a1a6b637b2dbd75e7e8204fac3db66e1e626cd4a268c9c8223eaf9009a59c553389e4488edbf905fd468d80ba1c2867991ea14682470c25c0ed452a3633852c7dc32da1dfc91a7578c674636df5f2d25e6e2abe6e876f8896cd2df9dfe5bb1a2fb9d1e7fdc8d53317865b645339d1838389f7336771fcfb1db0572e8f0bccfd0fd96f36b22515f92742ff7be5b2e682882b4043fc08bd6172f7affe238559f5a62bf61c7626cc12a516143bd647f582047c9eb5fe9f4f28b026be215a3646da5ffd1798def2bbe78caeb207e86771d61d60062055f72482124089251d7b84d7c8d68d76b3cd22c7cee49d711af68262771ba117f92925845e18baefcdcc7de831f5bd0fa05f028597a3253a3dba40e0ecef7d2e762cf12712bf6c084f6839b5b435801e42bb5ad9a893cba4cc9fc1eb957a7ab517dc2ec55568342747ebafc31052c17f2daf283827cd06cd040dda51f40ce6045e40699e14be926059b08fa34771a504e494718b412091989d240d5bf9c04e7a314d546d7e95a9ee404c20c3c0d031c632bd25d9c227cdfc044b7ee8e3f80ce1063e6a1d2703777272a9ae9c83cc2e9ef6a8ac1f566f5ba106f20a8fe31ff4f40a8f930a7a96fa3b99b4d721e6e92e6daf10e7075c40a201c2f0db130b49fa378d727b0a8f55e57cfaa456a949867e82b17a76773b97b48da890935ca555cdcfd5cb72edc30043a50ca67fa5037aec8ecca38ccdbe6ee45b56fabfe1cb2f85d6a212880be9d8a5902794bfd70205b5686ab9c85602067e931ef66d652a87d74033935df4a6a19869c8959ce39bb64ce665074dc02d88bb0ae44da1bc5c9f805880781b9f9ea615464ec86ae53ac34a019d1a155807d0466a79280722384e39b815016d31f3ee454249724ede13151f562807199bdf0c68b2921ad661451e2d38bab0cde9cbf81a9215dfca43e49aa0579c301db16eabeff490977e54651119d2d2d431a7db1f27f35e7c94c9ca3ecee216d7b45ff6ea5889b460db761a4d7d0297b6d0d64c67837a5f0954141f8ee0b7e6bd6022453b129565de1617052cb12048fc3e108f85c21198ba42dc0c907acb6da4f0b433b6c717c0eba017c509f60ea8294a34727252de707d2b507a95e3829ba5fa3bdb77c2c966a53baa4ab8ffd2e293711b8f9078e922b60044789a91a2fd87cbaba687641ff495110983d19cdc86e4b259cad0660447f067a908864b0013d0719eef498ae9a2e187f6fa8d2416f49d0fd409371f16d7603438f5fdba804a37910fa7b93d3cb65bb9b5784402f1fa7cfd48d36b6ea5df7f46f78b0e4a2459ee99f618633b7f9b1110d8189fd3c1e14bb8bec72d4e5039bf2313ddd0294fbf209ccb5c5323f9c2517554e312ceb22b8bc67ce08f8042f6d9ec41a4c4b38032cce888bde5e4bd9c532f94897e89f4d78a3e2f9099a8b5c7f74a5087de2c22855c6698885c43e4f2915c9c5baea5f459f69c536c3865eafcc627c61ecf8eac422204db71a173b2c507b6a13c95d3e56073a0fd6bf71eda0;
    localparam LBP_35 = 10000'h2351fec62423c0a4740754e300098ef78c6b18914fdc2a5966f59995f9b95d620644eb29c040bcaf1c7bc859bab6bdf3e4c9b5d6aac2d55eb8fff1cfcdf60ac2fa70640f1f7d70582b5e6863832fe45bc8a9c33c6e986f0f0e72a48878019ef5447d97cc205c8f435e04650e4127b92594f776637661c623162ce75120c89cf112338a8bab2154c892de9b5162afba2b27706ba626c46dcd81532b3ca10dea33aa0edc68e1703fe904ed63b922e8048f40183877935cab041a7241ec621552e4bb52a45f148edca5ffc067b393aaef173fa8a939b7d93ccc9a1c9b098cd45bbbb0a4c569765f6138ad72804597b1726c7b9628818a4a8f6eeb5bfddc3bd2f88a61284927b572895586c8a38a733147382a14cfa6b6cf1fea7d316bdb865b13ebd8d938a77107c9e962e242a88e7fa590a74ae7de5b5c47215a7d95f3b0853a6b1cd6c18959b603cd8a7d23187adc68a7d83e1261f818823e6098c410adc124965305348fc1da0e234d78d0432a0acba1fd8c2565f4c95653f41975a01bfd71648f4e932d7b48b05eb9e10e47614fef0978eadbf08a4b8b2d0f77fe324a9253391b3135513adae503c92c9c6b3fe9b0b281ec50030f83162fc2953f7e6c708bd34b2709107697ed1cd3ac7505bc871920682f97247ddbfb1ea99ca74790b4b2cf58f16335d9dec029625bfdcea5d7973a33e5aa37974418a7a1b8d8bc320732780d5a33a10d93ad19b48a28508f3e47764d7745adddcbbed2d1cbb88a411421374d18b3d233964ce7ba3df174fabeb06b988294ada0a5c9a781200b251815d04f1f94ab7a0272ee4f4251f10b19c3cf4379cc1570a866d80805e7892f6965607b08e77addb11db29f29d20b925ab745758c903878e9854cdd3928a1653b467dade90000302ef8e1e442e2c0cf3ca8d0cd1c3f4427225785250eb7678cf72b63388a0f0cc14b46874ff177a4728e885e631b275ab9475c8d26f27a3c2fe8cd06a0b2f4d8cd7699e0e51a1c96f699e077d3a9c8c64671218b73b06ea076b1bd0e1abb98a81f8c1bd2c892507867ce63712eee295b343f008c2d568567351866e4e953ca85708008538c393d086fce34e178718fbfaa1f12f18db7f2bdd831cb08255ba7f0ef8a9881e1a245393f7b77790d8dc329e9ea1c0333fc5f31f11f9cc969b5e524f5549096c92185363f64afde9ce31b097e0e289c67512f50191b39821b8f6a03f6d183e91b19f719bceb36760c219acacd28806098d3c3a98a338677d45bbb4431e5a6593a067be95635c3295473d65cc6654c9fbb3e971ca205c1f4ef1184913c8104c5f0be2ccfcc8c4be199b2252b1a5dcf75b9d1ff37b5130dde292bf5fe0b43d75f6de8af6ad6525f83dfd0027562eb848e81faa474fc97c6edca959d87d24475f4679d78dc1a1cc7670a94481ff954db4912b47dd12e0d91063adf63d14de044c7488176ce1eceaac5ac09bb1f5179fc52474b76efc9606faa390eccf6eda69cc757fc9658ebfb2c90096bd12d697822ed45082fb2a96ff07d15d8da87751ac3fcd4d4602dcf7f68ff0b9ee619db83fb79dbe6f5148e6acd76fd7b1e224a454557de97e719352c6ea70ee4b6bd484d7433dfc6e6e0ba8f427c5269dd89d3c24e33af9bf22c571379ecd38fa278f932bb81c15b44cdb651fd76dda1558dd06ac597131cccf993042e62c105963e2a748f01fd0b3287eb46ac0660a66dc1e57559b0c2743c9db457c4c21f75d7f8ac93daf540b26ab94737324832401;
    localparam LBP_36 = 10000'h954cfde12cce9bf353852b90bec421a58fe1a129b84bed4f638c4a7905fe789388a4b777da8100ef67d5d2002397dfc7f1868a31e9fa60c9d44a0ae6742d0cd0c886bf969d0a2a1527545fb73905efe17c6ad924314ab10945fd669da8b7b7a737dee961adda0e690a88e3670996318c7dd25bb00b65c34fc75bb2204e237613238112da5c370c431a5ad6b8b2c4ba2e97c9ac747c0adf988660eabe5b714ad1b55817fe339b6014713a98cd33d54e70b49538e0d02bb9c85f460492a9ff521205b3a1ff4a0bfc0552664723b5c6f5451553a710f17e84243580aeafbac62a45353b99d54733d5f10d068a9670f09a6a7ab7716330bcbc7e7f2e465413d38365d5fb706c187ad6150fbe6de5c241da0746b63ec8b2a2a6547a5dd2d98b3ada10c18f3633fc57dd9618507e988d14394fefc63a848d0ab953b814fddbb812d95036818e61263fad26187d9e2b958a9ee70de212351fc867b697b32fb94dcc937082f7db0c885c4e67c07761f842a2074f96b329153852fd5213d8d72e9bb2067dac3a02ada9ab3d4acca54cc1ef335eccc51808015f95eab0540af5b6398cbf0c252aa4cc3ff2561c3809125adbaa87e0bba82f8c8b6e5ca5d89ad76c7d018aa694a1529bfc6d58851c37e4b7f06bb16b0c56f82f9b70cf8310ce513308ed5b23fecccfd07eb77fb1e41552445b5d0db755aa6d0800b2a241d01bb993da7d6fe48d26ee77ebe22c245098b11fc74aa4c92d91a8f0119caba5828dbcb8250153ca6d8611a80951317ceaa607cb37bdb98cb6fcbd419f4d647d1bd11b1efd648dc6a79f46f22b99dadb3eaf580511445ba1e51815bc0df1ec2a280feb29a272e14a1261343b85aa73e962a25f0d0ab0c4c5a6e74f7ca510cbc20b9d3bedd0ae1e928f0409ceff5802c734fdb9ef902f7d0a4f413bed5f559014e3f8ca120999ec218f498bf28eaa4aa1131a198d14da823063d17d7f1d8184d1286ee9d501d6a37e09b946ebdc52ef78ac41367142153ec519eda7ca2a1f2f76a66494d1879c3f5d1aa6cc7580dc96644da07b839c20915f71e4232805d68b48da452bfb12044c23350305b36897329461bc780a006dc75fb66941a6c2616b0e84de527b20416b1049d9616391adcfaa4d667e511199ca0c0bc176fd25f9f7d6cfe9eb46ba73a8bb6877ca1cbc0649f6e97f03c9c1843b6cbe6888ef08abb60bc6faeed78bcf328ee8b69b902c90a945fcbfbc6ea0a483fa7283a1cfcd49db93afcdf405555eb04fb4c16e1f6cfccc92e8a33b62782ee7d968a17044558310dee8d386cd78bc03f080b81dc3c75280593b6fed89ecf09fb728544ee790992cef264eee48c3fa3721fec26fe1a3fb05355157e7b9437c96d521d659e8124c86dee201230445060c21cfbe6313bdfce23cfd9c3387d6520a8994278f89219b18e8cedebc0c7058805037d1afe9f9f6f99ce9c3da11197a9afc792bde5b1e53514f60d1770298dd096054ff3bbfb04441906c419669119721bdd53778257126f6eb1eddfa7a159703b32b2292fd34f51d1dff23b835bb5dc93870ff75d706e05ecabb968633942d1b9545cf5e0254e3da8a128d18ea712f14e909446b52bc4fc63f4f026b2dd1f8a4e0a9cd186a779b575995e3e7ef47dc61a58f122d3ecfc6610babe648c3b9735853c3196aa0239dbe4b5ba127fa24d7ccc03af3ee29b7d3fde56d380515f4d08af892a4e47b22e4dbfbdc4ea0a0d2aeea572bb7dbb28669c8378572742a4d0a73c414ae;
    localparam LBP_37 = 10000'h3d51bd100a7357b0745681625d9bbdb14e05e79a3fd68502c53f1fb86bc841c3dc16d32c33221fc6a1ea32a64f38c943df2aabdba694abc04378f9a065e85aa1f373a1dd1fbde824996d7c63395c28b63c220005f9a41b05118bb69d790dd93ddf11543aee9ac3142babf56f5511d2f889d94a4b7bf524164b9ab01a34bac13bd93b07d3130eab9a01ac95d7242e5e2a31d5906cd6623d7a3e8b347392450daa6c9ad5c9bce206d4de215ec384ab4ed73b946eadbd558d7f210c0328ee6854e07c0aa3c5ec188f1174379b52b1704984fb6b2c43f47c0b1355b9c289cf7ca4e8a99054ce7800b439ccaced27a110c4291d61194e80f9bcbbe029b6c49952a3cd9f0dfb71d9985fd94bdb3e45f6dd62f14db3c281ff84448876f60e7d81c327526d1516f83f68b0972bd92b28f32644db936dde71af383a37ec64bb53192e1180d3d187ba2843990d27d66c82595cd52d53263cc089c70e1d6f8559e8403209c155a757e3f607f3ee3a7e0904782b2087d598757b06c262a81513e793611276dd8a69bab26c2e548e59c14b8667714a72bee1405c5b3ed0fed0c0de74cfaa01d76ed2bb61685d1a4f8e4394f39f7f22865a46e3d69e54c27c72ec773741b50114eaea833d2001f9d57b265c33146196a8d70b1497923532a5f6beea5dccf32090accffe0516e604443df4975c5868fdb35a1ba495b93af7b4bc981def546f4540f3ef18c1aca3ceeaac570d75e1c104db74c116cd970a6802aee2f381a49b8cd82e2a4c007180b4bb62c58c3fdefc1ebc7cd6e2a33861f7dac38fe2474bf6383c0d4f9f676856ce473b9ab7b49e3cab8fad37e9d1c53eaa59e9fa27faf39bbb5a4c3977433a8e3cbe701b2fcb716a4ea85343e817e503ee3b693b26ebb8bd2b324a855fdabb7639173ef55dce6d6aef369282efaf1c1d004ac70d66a86ffed2c39389807d91f1b36f2995b3ecbe3d91117fc391bfd9880b4cd7816e47a6508462b91483637fb352c18ee29654901febc748ac6c881de37adef1f7eb781b23badd38502ddaf45e361aec6655996ce0f72ade26dfcfe4d680162459e50ea929d3bf717760b5114630d18f3b66e64ad71999c50c84c14efeaf442a9d153748920db46230247e9ac3038b414f593d203f9683f5bf10a9c698f50ff36f49950aa7f6ecb67f04f7f7bb9b00215831703629c010cd633f8fa7d6aae498ee1e354b68b27c402316dff6e3ccb81a531b640cc9f4ccfc5f4314b9ec1fb9ae836fe22c8334f6c5bd04708c6e3bd3f4c71fe609703bf649820aaee4102ed03e45e355d5f5f715689688404b507145a3fc651649ef574051e65d0ffee8020d2e24351fc2333c6e08368ca6be8edfdfe955b4d6be111066da4afbbe1f5beafa614c01131882aa1abf0c801d182909f6c8857233633a6c97b772669024f250ebde61c95668ab6e7c659067a5c27a5096f852dc37f3b1fe2dc28c3f023e3f4ff620b4a1c626130b273e38cf99b2f9fef2deb61883dd62b28e692931d64bd61830f91b46257e1f9336605b8616ef8b27a9232b2ad67cab42a5b2c5f5b809cb13f80042cb79c021c4c920dade360c76da311aa73efd103e7b0663336065de70081656edc828e9f525ebac504a06a76c38522de799521cdfe413aaf79990cf2212488518156f4bf06d0b9b7468910417468148f05d4ba78660991abdc4f55e88257545f80ee11eac819882d62a6831e14296547e87e04431994127dd7447415610ff3a77f605302da3c4aab7;
    localparam LBP_38 = 10000'hf770c0cc80f1adb5e5e659dcec215549883aba27ced40f2134947d4ecb45d222f53008a7146b1ac5c5b0e4f8f6dd09ccbaa5c8b7ae0d1e92010af846469067b52dfd71fbac6d8bfaf099b488070b2d4b715ede9671ca1398577d74bfe3eb8f7e3e01039e5139becc3e27b41f9140478e1f9b0df9b0c2d24d9c322e1e69f5f02f8a32ec22a88052d9cb426e30dd43f810f36ee1f7c53f4f465f4468ceef15af270bfb5f0aa91d1484388f850cfa19cc788dbba9562a476a65340d711bb09b5be3fd290ece29eb49f1797602c53442b0b673bb76312777b31d4cbcf414e159740a350aa1b34d9482351cc6dc46ce4a7112f58915c49b51072a782a71cafa7969044e10e70a4afaae2b83f4d44959e94777ff3e431ef5c51e3fa0309cedc5c3cb55bbb3757d43e36408aebe12fe4538073cc135781f42eb71613bac15fa9ff90463c53fa1c689cd63426ce4fe62a7d3b71163f47df6eda06a0eb9579be5526bab41115f9df3049a88e408f80d61b1b77fc923e192a361bdd3111bb602860445143f2b440104bf3470ee85bddff4a35531fd3f0a9be17471e68dec3ca6edda13cec72b9ed91166d74ecfd1be3e98693f60e9a91a435594c77737f4f6a50a165a4b400188c657255b663f1a72e9e6fcedad92b1316a8ab4284307051e5cabca6fcd8d4a64d95b3192edd83ab6a261c8f4b907dbbf38a3544996e2200a26f3db99c14e3597a39db38be7bb71e3ce843d956d3ac8e8bca2adc7d24017b9718093fcc2986ee464236911e6a096472a6697094a0832b2f5a709eee281e6ed2be69b2766a0c67565efc7a66c7d71343d1e1679df0d44e3adc44f49e4e95a7438532e27801f8303cc3bae2eebe8248fe75dea2f375078fba3bca5d634f2a53dc9147a417952fe834b08a93d9d008b3f188d9a9b7f64c4b49b14d1a664b7c192c65a3da1f588cd8fd2161f7906551a051ed2624f3bc737ad0458b8a886b2cd11db607dbc9744bfe4dc60667891b743f21da04e9c5a40fe8a002a58e89b57062dc5fe638563e6ca0e538cdb086a4f3726d3fe690cfc01884be3dd487e901cb054c74d6a487e86aecb7258fc88d1935a257f90b927100f1c966c822c53ca4e6b37b070940e4d0424d8d955ae667a3f2e964c15b967ab263bc8f41dfe20cf90bf103b66782cb13d93c35a042b4493c6da947bbdae34bf03c8a0ca23e7701358b4b84251db1fc3d1fa41bdfb7bac972bd988b82787281772bfc0ab711c5e0049562521c576d488d24ccbe2304cb761bdc9536d8893784d0fa1abe077ec9762c067c4543ab0af340d3eb2a5d90a3c66ffa5a320dc1b65315e64514554db39cbd62fd92bd41905b676c1b09efbb841db251fb0a1ec97fea19fcbdb6dd62e658ddacf1e7804afb35d70128635afca40cc21612928a9adaa0fd53b3fc174ad0025f7f50ae06c679fe91762d7ed9730941ebdba3327321381c801c8eedc9d4ccfbed823df2af94d772a37e04af238e998031a15247eb7dd370419cc4691f89e9f9862e192a74508753d3e56b3ee59466b0b375b8645737f65e57b01b37c20f478b82f2705cef3cff9947dad4e2248b87fe82db5d358bad001a088de4391346a408e7fe2368b8a90e479b1e5d0ad156080681f75f6fb81993acf331ce923086815e6f494d08282695adb66837c4acb813a1c2cf017476677a5ad2230e2af2a9bd8b02a07cbda2d164e28e9154454f9c09d649e253598ab07c99dffd813de00164903d0873b1f490d2038dbfb5a;
    localparam LBP_39 = 10000'h155fa8c1e0447b21ac7c49b607cab186999a0eed0f3f85cc58a95517bcf44dffd95d284a004507f8f6c260037eb421d3d42124e06574b3ad67f62733cb2c1523ca8d2c9132eaaed89ce5a5df07b17f92bea262e0aff3672149f8f4462900b46f1c1d17ca94fb6280acf3d2ecebd943bee40b1a35ebd03e8257bf72594e324514b19769e93622b125e581533d8d5c3307b5be3afcf5dcb43b184385ae16a6742c34b9544eb8573fe21f689d7f5218cb04353cd1ad03ff614b48bef98088368f534457ec0444a1180f1a2c01d053462ef5dde860d5b16034ca7f73ce60c69e3c5f9d33e7441014a402911ce8e74ff186e96530719b8efbe6cc3b8d60695a35805deeebe40ed96886080293dff832955e793832d1186b5b0e582b857bfc792dcf47ead1ed6244dfbe9a6ed15227d8872e168e7e37490e41136d1aac7980177ae635aff266651d139b92da86904849ae34517cd3771793eec6beb72cd4359db12457b159af6c75ca0ad95a7b3077123fca88da53ac6f4f9b9501b170b86a60ae28aa311400e7f8b98ff9b82f7c938f5597340bb65c338ee99a86060b334367e71ccc3845c0b1aa8769881dea16a5a2fcfb02dbb11dda46641a365e547d2c95474c3ae47332cc0c184f9e8a4c98e06c3eedfc83738be5abd2f9ca8f67a338f3f0e89320efcb407a614b6980e0372ae98278d93bb5044d18776cd72b262d45a21f5a74b641f7c44e195eeaf415dc9632f03396e30ea9fe8b860d0528878f75b67658812fe36542e47b8e37bc8b76fcfc17ce77f725752b8fe815d255b316def80c59d3f919eed92e3152d618f12227e4c1e54d154b9149c5b69df3a7aac14c44eef2f0a481df0e6e330d8df51adbc07003e9dd82959f5d4c5ff368fd5eea9da421c031a1b3158b584458161d7b0b596e3b00913ccaf312abc7ca9accaab9482e07a368bb7855b3514b39c895bd9ffa75d291fee4a39ddc27e5870923d58b36e881625d483c7fd6706ad27349b8cc02654384bbefbf33e826d00fdbaf1214a30b1f30236b874e9a834232321111060f5d7b0719baa5323ca3c1238211dec00e305989e2c1194674ac373a005ee673e7573a4e9f86014d301c27570f31fb61754ad9ecf7b225322d3960e1ae6005c03ca7e0ebc59d100f80e6c8528b5ca6db941151a5c197822b828f964ff465b3b5f3bb25bac3023840ff134373c6d83ac61b32a6934dbce1476c700257defda3de943b66f6579fe45eb1d95df0491202ba59d672ca68c4bef8b71ba30478df0a5623a68cd7aebcfd3dae91a136da54f263efa764135504b19fa8e2c7d6a6836399abee5c7be1a942ec5ed4dabccc725d4044a5ec4f5c506800124f0add08b2a73ce98825962c59aafab7049e3910cb102926624454d6f12ca4967bb6ba3259ab6adc196cbc6d696b029fa95c134c1ee7162753432cec6e686f3e628796a91cfeb95bbda2ee212226056914d32c0d0b413ec9b2ae0f57333108d55753d6669f4b493d0bc3977635ebbe7666f215e8e26f86544bbddbbc4c01722656aba66bc64430e24cfd927f18b260813ce7bea92714693e7140274313e395a6e4f16a87f485e9cb0e41560351813a1560c96e3a5974bf47baeb461b6c5145342fd2ec075eba4370200c69f6218378e7f667975ccdef9ef1e1805767cfea04eef4ef35bb2300b766a5656ec83cdfe6224fdf7c0182dfe6c2f9fd670f03486b1ebcfe9ed3a8ce7d205480675e6ae61ff503dbb434843f4fa20bdc185331f2;
    localparam LBP_40 = 10000'h11e457c464e63700d5596405220709755bc0e06e6bfd5893c85f72c8172855564fbbafb20ce268da9f6af7580211b17ba480a81aca6fe694bdb6c974a7b48b8160ec2a9f4fd1d549a252b65aa1c71ba638b82cdee3f9a1d600355d99966980f022f37a6731675eacdd9385c5d5e4b832bdaa1968daca0cffd1da6f3096673f6232007a8d543a39df5a2cd3125cec477650c5f7426fd9cd69d8ebda4c1bd8b431f5dcea99206b4e5576bd96f064b7c2602aebec0a07479cf908b6849736c02f4337a434dab2a44601f74ffa301ffde4e6fa975263253cbe2c9c18e9302ad3f5672fd0801ce27b7b9f444fedd7f33aa114b87ca32fe503bb2dc0a1d8f20ba8dbdf249b326d40587d4007401e2c5ca26c58d8f789ba298fb703561b4f4d38d89204bae9ce9cdabffd7000e379750ae77d6a08ef6f70421d80813b039f458d3d2d03eda49f243a34408dd9726e56a36c13edd6448e211dbf28b6575f4fccb1f6573450701b8e0f3e5054b3806dd25805effe8f97022724796d82862e5746562a93667d3bab731d4b55aceeeb0585d76627bf973942f331f7e0e99e5c6687ed9a6d9f165102b54d41cc0b9248a37a1b404434d0a888c468e468abcc11cf742c52fcdcdf2c8a728a7f62d6a0e75e9307e90c2c2ed3324e0dbaa0f0b7425a18a5609e5df126d246dd3e3c19c809a20675196887879a3535871812bfc98330a13527d3a3f724ed98d1f13a0353c8f10353b73e60fefcc7aa35881bb9d3748cbbcedd3ec9dc4b868b652df678fd7c4a3fe5bb191c8edbf308e6073f108d291f235f053424387e27ba267ebea5d0ef73e958ef2f86e77a947714b2f0216b5767a0bcb9ef9aba45e5d5404ac9d826a2f80f8553ebb7e10a2bb43866308d5ecebd4d0cab3992dc1d289d94ec2078cdd3a58505bca6dc40c2553355dc220b622245fad62d4c166c0706ec83185ec25222a75163c3ec46fcf80260f5640d221ab57ca780b70daabf6dc3d7b00606dc87d595d0d4e3bfe5716285a9bbfa7ea11377a3144ea26a689e254900160a5227137707987bdfe6f84d9a01d90be7f38c6d3e7bc413c3650e8610705f04971ec6c2510d12c57b35d842e71598e90a64b3707b8c90fc7364a24f80157e9260021f4e349a9c6d3d9bfa9d46dd8ec74b24343e28cb75872ce1a40327fddd0075a4ac5983a88258ede78fd75a48a41c998931f862fe7b2de018fbe5c19c053fe417faaa33cbd58c43d8a1716d97fab41c498996235346edbcd3a41effdb8a6ead966c1d55435fe2efe84986865c278b07b3a9b1cdf8d1498be22df5b410164ede7819cdfd8df37fe12db258d83d7b37fbd36bcf22fe47d0349aa1d02f45d4ddd249cbf40fbaabbc9ff052b931e08635a1fe74510fdbecaf63699238696981162458c840e68c0f8242f06220594eae7b3302037c7dcffe84eadd8e41f14fffc05bc3d4bd9e64e9c8648fae2572cacf09a9182d61293947961bba2625bceb0122887d2c8422ef7341636a89ac26639bb7c891c75831f61ae7fa86781cde0fcef3b327f13ef80f81faa07dc71c9ce2486b1806d14a2e09fcf3f054dba8497a5253fc95b0172ad6eb55317501a6ea7c92c0b5b7327f53a9725f49a0959cd88726ce83f45678ddf85d218d4384dab271c1c1bf60a71d9a25ce4753d69cd552fdd67d3d735a5e702d424391b90aba80c80c5e651a396b9d7501f445f76971a9d150819ee055f92514409363b79ee58997b230330c0a4045594d46503fdbdcd4;
    localparam LBP_41 = 10000'h16463b6b418f87016edfe4d0325456b4d6c0b29f8ad93941d4d65d2e427be3736a170cd665a0d706af3cb2dba4e3ef1ad11dfeb8d5b9c74d4978a55f17b2bb9b5f1a94467cba91e8830e3ae44901f813bb8a226b8252de44d5a484c081f3e9c1527dbecbea2caca7cec94d8fadbd554ca6937cf556d2e1ef21c9031fe5b6f99ff2efae1d6cf6f34cfaf1f0d5653a302c7b58e00924a9e05aa7e4ed17c41f7aaeb38e53c7372be972eb060e326b622f3bd4b614e162d25faedac7fadc3bc6c5b22f49bc14d1d46b335df4579e9e47d94945c429b353ff53d40c7f756927f696823bcf88e0c6fb1ea11a9c10722349549477581dd9e49f4b335857c3e2d9066b319964d6bd37c2766be4b918a579028a948cdf841185af0671df979dd9058fe6c447e04ef571f2c74057f44b5c786add86f184e7d4b1bb1a401828008b2ee4a0f3c966626e75f5e266ff2330a7e68259e4cfc2f6245d5742a03225f932fb83d25f60ced17d8993c0c1d3418631cf89ba987f6b0a13adf3a9316b4c451b532a145a62999451a23265cedf91b74e61adc07d061419675a763ed00c42d4ca0fef7e020a3af1400f87ee15a1434f9ed5cdaa880fceb4e4d1028ccc8b4f4831786acccd215b333275d9ee88f1b40f5be7770a89b4e890b93e0fbed8ed7f87150472062c62b72a7754c079851d6db5e778e047d9126131e55e6f716411513c63b0f493f78202008efc1ec487052f58130a7a59c4fb63371fda9fa3d7ed6fc01aeeeb59cae2aed475a0e5d4b6eca39066e51598aef84bb4006118b8af52d21434641cfb3e4d631a5a1e81ccb62576f6dc71a28a400128b238961f9915722db413cba496d76834e2b046d891efc2362df97f9007787a331d2cdef1138adea51fd64fe08915490c1a62290493e861cac5768ae2edb5b9d4eb8edf7d08383c032ee1825bc6a2acbb7b730b92671e06b03453a3be4aa12cd4ac0d97d009c59e081cac40735d3d6b584349881fa102aa9621a1cfac310915c77fcc49220e6afe293561075fc3d847afe6bae1a000a32455dead4bdb5cadb45f8812bb30d825281fccb0a2721a41e76e6c95ff57c3f44c9c426cfd1471db63f9b0c74d142d0e7eb46a8af159affa4a82f67c5039036c9c1aabeafabfe06853d84ecd09846df133c1219207f1ad7bacab1a7c9decb642d7e568a24286e42cfb49f0815e0ea4ed76a2e51698c425a62b47b28e1e325702d080be1a00909b9428f57a4dff906d19aac0e633daee902dc3495b942167a3400ba103d33990a25e1509fc2444f8db8d9773ef0c39793e3cf8597fca107d761c075e935c08a113513a41c34de57cae3b137f1e2d943b0c7dd5ff358f6ec2ff2dd8a1776ebffab8ee4c2cf1a5f3eeed9f14cddd563e323487ceaa70a8662ccdfb237ba28e20432141c182efe7bcaf5faab90400ecb0d29f1c948e4d9b07905a42791e6bc65d51e7f9dc638b961237ff9d7805d356335ae4a8e2505ba986369542e172a1c521fef2ec7f78e9e881a65aeaacca6b844968833ce4dfdf7e0d911a53d165582608e4719a6b372ed3807b2117c4bbad10fa95278d32c90aa2333d37d002f8496a85a67b3c43fa51eca3949c4aa015ef5810a9526a4cf093c8d75bf5dfcc1157c6fc266bd80a96e32d4fc7ce3f0d9730482987481e3e61097d7cc97d0cf40e248fcd53f262d60be8551df9907619ea49445826d51a17fd793f3b7501739ca452b4546b692479e5db36779c5d0409250f81e888bfa5b503;
    localparam LBP_42 = 10000'h487eec44211269a319d7b94d41bc25424ea199e18b8eba8df17329a9843ef8c8ed546e902b486a7daba9c2bb0202c1a4422387792776551917371fb01045ced226f348e2f724eb585a0d29dc03f4e78ff567354ad59dbf8d53121c9a2bcf700993a99df0fa94b9853f1c86d7b4dab34ffe5fe810fa4e7b3945ceea00019f1960bb26c58530eba6f1f4a48d8f2bf337e7ab2f7d522eb14f7273e9f3c314e3fdace809aac95be78531f8b011be385b3072e4d7aefd556f39b195a9b1262f25cf28fcf0959402a077182df7eac68333a4534a9e8e1dd8a0a9f1e6a7d6245ba83422e68c0ca2c96daa031b8a084abb4098c08bda1a5ff3b8f0455fcf68726d87f66a931b3f56a12fb06008a7c107d6c1953cca208bf14c321ee31ac514dc841ad9c39f2607462494a3fa2c678fda511f52d836c0872661af7bf13590b96ea84631d411f2e319d6c647789489fe72c8c932d3e8d29712e36fd677e1fc4fa07a5dc9800def31560985ab6b46f6f982ab4f56798091db03669918bf926b706904b1d68144461e26b41de82d62e42cb9e2ee4089c3371cc28ac32363f48e112db04740e830d56e69bf7e750625ecb11e7c419348caa82299431680527bd4e79cbf7ef002872f9c5086a1df67ba9f09bbfdbc09de9977d8716c6cc171e5b63d69a71ca00609c85042878c0deaa06c89bf1986a25c09e092f7dcb43d4dec783957a38af73edaaceb4260bcaff107da2593daa136c84f03b7846fa7dd1f66612204ca2b4cd6cb9d26692d40ab8dda2ed8d62abc6f1d62558668d95b7ba5808d1b038881b4dd0cdca3f7bc6f081279db2ee9ddc2d05ecd834320cdb9b7572051fb851644785bb1a9243bcc29bcdde0961450d8c69aff9f6c4fdd25bc1e148e5181af08b1ad83cbaa54f18911be919162c80d97bc1f4532ed97c93ba736a3af041f60bf5802f2c650b365e1daf53ef958799ecfb1542686f9745fc458494c22e61f5309af6c900f017bf1ed04434afa47b4aecb45360b9a372922c74e964f641d6ed29e02fc170be69a8204e8bcf1dd4516c92b2c2d05aefe5f31ac63d6b84c18b9573b673041ae2e1c783eaf96d7ec6da1834cf3022f3797add8617337b4e80c29c13c86ed9adc3500ce624df4eacbb299e734f5d5cf29df33c399b06192631e76129f754f4f99cdc3eac73f75a4dd3b8a6977e03591c2ec7f7d76e14179585f1622e5f8df5828a84e0a61ea7834fa0ff911d464613808cf37f9d00a58d089420046f3670124df61545c3ab7ff4dc8d1895df3f562eea84c381b345b0c8063d54bc9028ef3bf7a44af65907bd4ccb7cbe3563723139808b90f2f967ef439baf47f18102cad37326e6f2a61563a471172f86cf3f73a28c50b9e4d63263bf2917cbe1b03d04d8d36d054a68484bd8542f023ff74179295b2547c36c83edae2994cbd51ff1fb4fd99c4afd72ccfb1eb662c203651abd2c04d1c9905e77e615506a8dc9e9d12a5ad887dbce06549f4e10fe6f6460bee939eb989db1c370c97db77c261b4fa7b9aa9cda6bb548871376bd88f26a7e55e90379fa4d38221072ce23890eb17a5b4afc0e35ff7923a2030ae106710e05d8b28cdcf4e8c944ffc737a9e15abe32966b09dacecad8cfc10ccc94a3d98891e4ed019a42b533d58be1eeef0a556c8febbd8f8a410ea9c44090901129c8b76f26d766c8870caf8205c20fe333c3f8495f3afba5d80aa35ea4883811a545f9cb6d4b00652e9771e7747498a8763e6e75c1277272656;
    localparam LBP_43 = 10000'h8aacebf1941488a7869108bd65d63203c610244aaad81bb7bf0cd5c2d64dae2e7961bbc1760fed42205b57ff5aec700bd52ebc3fb6e23ca58282f54f6bbd6d26abcb3b6fd2e2d922de6c0311cb2fadf1e28806926b6b821061dd62d19651533216f58bdb05dce1bc64e6aaf66e3e158ffbd75c9cec3ad38c2091c835be168bfbd86933e3a6f0d64ef31afdf69466ce2612fcac95a9bbccb26ab28abadc7a88a2f60fcec144f71fa82362eb8d87ecfd80faa2377f6ec36ec45f925d487e0754e1d95072c1b3be5f14c2945cc9e4316b62d528ccf1f73f48bd37488e3944221199460cf19023ace570ace62d4c8f87caab4d694f21c2e9d2023a7706629bd4b8b1769a87e8c00de7784d53509b4a917de923146bb9383be6d30b732fc5f70d3cea7526316e0f760b53ffd0fcf4ed400c241832bdc469f0a44b6d1e8cc9052ac6559f92be9d95bf2b79f898f56c581eaac82f8b4fdd3cf521aa17639733ab47354f7046d526dd10356f1a787887c898c3c85bf40ef2156d2eed2846ebc1c1da9b0623e602eaace7915a75a512b6ffa1c4a880de8db3d84b189cce4c6d1caf9ac974a94eb3a381665c0e77ba71a8b45403f5aaa46807d6ba5f83c4a99bb26648ea5a90b51dc85f5a7f268ca5debc1f80f7c6676aaf061f15c06e103b58efa992f5f985ac02ff1c41a8c89a202bc838b31d841980ce82a85412c00b2a523924ea9fbbbdd992659f46a69729a7c4c34cde26901e62ac6a550be0c913877831b3ee596721aae690d8104887231c11d58daf5a0d65e8f4c4ceda65a6eac8a948d7e8c8cc87ece8dac4637d90c0c8221bd0e842e31e86decee62fc54d3934c52c7f65fe6a3d7fed713b0aef5869d78f3eda897fb1344decb799fe99b2c323863c257c03a3581e13a8803add8db7e5731a23cf19ff312b4014855011f81ef29e4d2c1c27c2651fea484a165dd92b193e0e820463c44cbb1d6a9f5208ecc755c22ce392b9a55dc0f856b061590574fffb75ac6a40b6cf92b745f82c04c9e7c69261d6b441f62b79de4a89de5f6a6ffbdcf30d6231ec4b719de7659bec884cfa013194601101c7b6e671467750712de8bf9bd9d2ee57fb794803caf073e0441802d20a43deda0746f84f035d8fdf9f03673ad480894fead70688cedb840a6badf94b264bfcc6eddeeab4f7e7eeb7a1dc9407ba16b2f9e824e8caa7df1d2cf280670a20553a9fb4d16cbcd969b0cec12df02a39b60b231f4153083b40e929c138240aeed3efc44d45b4a7e2f4c5cc6ef290f2d9140cefec0e8820d865dab15084253a8ea290944dd4f134daaba37b3aae09e322903d00ea416db7d2b6e9923507d15f09dee4f489f11fe10245c36c57edeac2b99576f73065fc5cc416f69f662a557ba79c44fb1a00f07ff90500a7f5bde503065fb8d23f1c2dbbeaa3dc03fce31bc7a7e8b60f18436d4f0bce09f35c22f27ec18f08ccb576815d5b7480f8889403e395492f2111f33770725cc722cfc37726113e5ff1abb811ce83168ca067c018f872d82d41aa82191412014c0285edf9f10042c3a4c23caa3d08835bae15f4f01197d60e5f06c3b284f7d9875f09195a96d9e01c32ab4aecfda45cdb29b3bebf2ef194330966e9858fcd3aaf622923510f8e9f279c6ac1325b7b7810d0b5f489a4d385649f4654992d72b6dfaeaaf9e86bae4f06ce125a46f2b0b9233655661a342475854df8b119bcd7740e2035ac32b7931377c2dd1236f1bdd04e9ec1b11c80b443f7c8dd40;
    localparam LBP_44 = 10000'h3c9996ee649e8b98256244ed5f09b4583eb6142b53a66e44204f710b00ee5e2f3c2273c3a5148069384d56b6adefb9c49d3c61c6b269eb78993a7ab4b83aeae7dba4aec83c65b0d9caf505b75bd286a0d30bddbb5a622b420f11e0564f31f11c28493de3c7350f8bd3f2e58463a8a3f390f1114c09c48d979839aa9692cc67d013752e234e279b4d75a9e08fb9d20d11dc3f66fc0d0b57e1108f64e4ceb6698b4a99f54cacb7c3a55f2f662ce075e0f7cf30cb19b31c0a1665e26490a5dab7e5d65f1dab9f57ef6d5da8059b31c792646c777d8d942ae97cba66286c16ca94859ecc4f90937f2768d40ed040c7d289d4e87ad535b22930f7717131ec74a6d6fab5bd5483a738ce21fb5f82e2c399051a3cd05adf5d25789254afb15ad1b24a7dd53da430a90b8bf6fa94ff8419881b39fca481a0ddfa2806c42956303ee6795b14f30c1f78badf2cbce7a786da7bac18fb64cb650680749e1da1fd9860eabae2ecaf951835bc9c3c65b8912734fb1b4ec7289a02281df1a284d15f1450cdba1ff8d929046617d034577141aeb5fbaf09552088265e5e0a6f3cbba3ef0fb016c0f72ee28c244a2235c79050c2f1f970540c088be131709ec812fcfbc0d00b5b1f519e4a169ade275db3fdcc05700c1a99b852b47379357efe66b4835f1b5e214c8a68bf6656854f8b279b153b86bb3a8d258ba8bd8f6b920412c07d774f12482d94a815394f65bc2bfbbcfac69e51a52a41601ad997f94583efb55a53539413a03fed10acf038f0e75bfdcf3c93a55b92921a593521539c7aa4acc2f9dbe6d3d86b632bcb4203c696696046e06c5abba45a91e104c70c49887d570cad9ce0d807419cd5312a244bf6a30fa7b0cfaa38ab560e97f78a5cdb74454015f821893ea0b58210b9b2ad8717bdd0b1091ebed02eaf2f5cec0a4fe10b62fdb68d0f0b83b93ed04175bdc503c1d4fdae89c4dd7dde4468d8cb77b4078a4d83b24bc91dc6055be528ebd561354ea943176c1a7026881d4827a498d9e86e2772664bcbbee1b3a9fc7aa274061642b6081c121d282685895991fd4d0b041e484e690ecc9113238caf97e5f154c2584d878a65ab8bebbd20f392b40afc347b32fab9243f1b4dfd4ff754a897b3201341ce7539258e40e5c9c271972b4da2a6861c8ef3e54b72f04fec7d51a2325c98dbcb206139a83e93468cc6e1697271d0be309e837cb0ee4b1b241b5cbafb3cdfa7cc4fa6bbf140734c6570df6d287cba2736668083114904ec242c399a104f958af556bc0877f6afc1b6ea7fe10b2c3b3fefd4a82b9d972d038aeaa18eb7e05531fbe8b01dabd4dfce540051a8b9badc83cefd591dbf61ebe90a6ad30aa78b0d49d51e273ffa7e9b6724db0c569518a7d0eca573c91ce5f2b4692738233d4b4035312e48bb1cab2100988179bf32b2f707d2fde3abfb08c913a3670424e57da3d192da837e0b036685c8deb54825ec71caf2ec0094a0e83df5bed22b6dbde704469909a48193a78415911f60507d9f1ccee37ae6aa45c12d985d067269c1624553b17484c8a785716d07b4c6b616a5f6f7f74626a52060b3f8fdd77d81801c31959ef94b0a0bfd66fa02848a3300c44bcafdb4bf9161e276e8e7fe9aaefc29a1334e991b1d032e7a6f5f3cafa5fe17be266dc6e8829fa17e91065a2b0b2ca6efebd9ab9b0dd628d4029cd4ea1a93021d9f6168c450d96d73faffbc68c8355f23ddbc284b716c0f777b9cf19107abf58ded3d456bb538516dd013;
    localparam LBP_45 = 10000'hc061c3d8ec92ac99a1aed482cae36e0bf90a621390bc5836d8700875c9867b096141b4bb1f80f482413c5c71f3e27e894a5de4469a1c0662c1556db450f02edf2fcde44fb4b47da58b4cc10d3c56e585145bb21434bbf678d52553163ac5f1ae0d2a8accb83291f86a7681ca61f9fd8a7b998aa5e12b1277f1106d34d63244a8af7d19d0b9389ce62f3445a21a7b8d6b32bfb3d3c39fd849705a16dd825365f7184b6bcb58d27cc12d1c1c604cdafd0866380e149d570498d012148a8250080324b23fbba883bd43051436446cc2e76452deca39e89d77b65c63156a3401fd5602c515eb2891a69c90fc3423eb4b16f535045a37e3cfb6ae517a39e1842711ff3bbabe9cb2aa0375c73fbaf643f143c6b6c166b4723804b1df47a782872a64613c5be9e25d1b5d2159ff6c5fc076d8b9cf67f3d8eaccf0596ac190e32cac461089b7bbecca26ffcc6efecc52d2516ef7373d68ece4c928dce8e0a8a423334c153a04e07cbedf55769e83ad08a251ece5c934caf5fe7d63745ce80351e92a7ce1e026e03cf29b31bec4bdf52f358118bc88bbdfa38df8cf53b3fa52231ca24f37ba98ec2c4efcb44b89bf05c85feb22ec773f5fb44623bd0e32df894d5f90aa96baa2571879b6efc32b58e4245b310cf6566b4f2a075bf36ed07ae7e99fc59fee22901193baf9f92fa81a5523fccd912274758f41be9d28aeaec572530d8fa323963dc195926321b81104deb10b11127cd06c865e201e009a9a7ada6aa3966a72c0a716f69f2d3b762fb47fa1cb2fb3b012ee6f1fdbffb06c72efebef24de898ed1f3297989d0ab6bdda90e2fd9df76b5edc393fb71f389a440e8c05f920aa1ba67d3a8141b91133c4a4b16fe15aaaea4402308b8871cd78144ac845d8e02545d1fd20864642f74dddb14a4a99802fbdd73b188a4589fc3991f3fff88f3342b7127ca04869dea9e3ea639c36a452892f5bf904cd0c4bb91c15a58eca285d2e1d25deb4a26442aac0ba42ab73752693f606d7fc43f2eecef97f0aae4316ba7c254c21a353476f4d57d524eb964ed8e09dfb56d1264059291f1f97ecf73450e862c723c746d7306ea12b2ab6592a0c2979751bd7319cad7e92124cfb38192c6c674c20bf6ac44c91a7f24f6a7e20ea34c727d08d0edb38ee979929213f8da050472d47703ea7b01d6bc972bbff6ead135ec5cfd05456baae4f74e2cfee55b84ad10ed42b29a970beb9a63355ef9583fbf44267047b8425db34a4579e17af843c6b001c5f4cffc7f7e064fa8d0635dfd68d9336d7a8bc759cca1e2219ae6caa0161028681ab16f6989c8d670f0aff769dd404ac27485eb42937809311df1ff2d3a42f64833f7e38211923dcdae570a245f52d612370e095da2a796f5b4f62958ef62fac4e8e8f1c0647bdef6af15255904c762496072efe0d176a1bb12b091949a95200495e3a4059ac0f8ea080161850e4ebc8ec0ba93ead072404eaf151777a8568485ae3bd8593096f827797d858d8c547947366446f88c123ba83f7cd0f3a378ee03ba1a8f95d449d0d30ff1ea5f18f9d10e0b717374eb370da59d95721288ca473d4914b407a7b168a1893e3bfe5bc07940d3bb45a7ad604ae1670ba0be3a4f7062b55dce9a157dff4c36779c8090cddd45e28c1db835d10e066413b22ce2348a0aebd07c559d0488c7f79e134ed1595ba80fd6b4ff13d3bb722f503a284b1e09f059634ddb0994f86b3466ba5245d013a38995b323a87374661aa9a01308dcf04b;
    localparam LBP_46 = 10000'hc3346c8e5d30586c9e48e22f01e0c1538afdf62e5942514c58e0cbfcd0168a2c9fb9be2e5b1a130f8c338d98a50358d12c6eaf3c7ef5302920235448e3b99c0ac813198ae0b56259e2c950375c0895bb87d02d01349b23bb81a4b26a74a606f8ad0c8e9b4b1b446ab5b2fd376132f31e8888d45aab9f4ddc9b5cc433cd5c3d371dc8fac5a951d406f0557dea809bc90b21469b09ae74dde395600eb733784329bad656bd78ca8554d059a124209cbba9ac3cd04045cbd5d6b7ed127f2de18cdb1b37aa8b2cc6ad129880c7d34ce4f63a76f2cf5aea4370bdf65d8c40ccf61ae868bc17a1a14c456a9ea5c2fc4fbed82b41dfef0d73e994f4df4d7b10f27fd8f484a9aa8fa48104fc060c714261a8bbdbb5598a60d6c2c810f48d3b231f4d42816273bdc1700962aacb256371e2dc289ff8279728098cbf6b472671bcdfbdc2ab72e504e52a786b6d4ae2399aace072538d222a0827585e9d419544be62e8d802891d18b94739fb2668934dab953bc0be8cdcd9dd3d9f5a45dd6a6088f1e9bec5a83338232468076088c324691f49f8d2d5a40e65f4544fcef1cd0ca2f026a63b15c3fcdc60fae42683fcb2269cf10096ffc5cc910d365f8f79557b805ff3141868d45259182c974e657f6d8b97e9df956149ab2aaf624535632d163888dbdb9ebdf026fc35e8f5e8b0a64a4dadc37dd1809e5167fea0daf1db272bc52a855e6cc3a5fab7fecf705bdb2a0bd327086e7b123fcfe67b15a3bc6cb9b6da23b870b78191af50671b24396cee762d2e1ad10285e21da800d1a6bbf20cd3f2bbf7971f21e694adb6e32fafc2610b978d618d898ab4cdfdb24815485a3109b3e3e2dc898b3e799e8dbff0d8fb893d8267158eaa0505152e821be4416893ca4a8a32913cc9b60a5ee6f65daf9c7e8d9fbe8bab448ef2ef90d43e7d8f0913ae58cbd8a717abffb133afdefaeb9fd1e35508f8962567eac0606516a47e514a294bc2ab7929c54624771bebef344b74a580fd1691ee5395de4946ce0eb4fca89b30982064699b0e40301216d88d35414f3495b9b8d9ab314102460b2b56995dfb0e649f356dc1d54b81f6099dd75437b82c416946669a84a7e7c7808e2688708716025d73cc6b8a755f440b5ea8d3a4b4ba5a99ce7ebd3089b3de228e1cd72854ed4322fe930c4951fd6283b7672530d1c8c6d3670d2240e15828b9f9fa48786d0bc7bf97fcdefd0dadfe6c5f02e79e250c966c1368852be65fbe422fc8d8cd295b3fd038a11a07800f573bda2e2e5a8cb00365c918b747e8ab579e48cbfec39707f8fe0588d3089b9955f0d9dff179bee93562ef97a671ab49dbc273c2528dfef672bd651868fd7b17b027b5fbb41abf54d56693d354bcb9c605b85641f245db462302b09445613c2daa2af6fd25e8ce95430dcbf8c4d3b713edb52f60a229727612218ec999c213b5a97b5b318584647954fec5396acf1e36ed6177013b9fa1e7f8d4769996baca2fb5cbc11d68c55c59fddd8093f47dedf6047bdc7850d0c87cfb687013505bca3cfc161ddb0c316d27d05f04980628e76049ff868db6812c30c3084067d803705c18e5ab2270ea64381b21e792b3ef178f59075624b7bb190e122d77ca9691429a11cf43175474bdb5a600dace6245d92dfeba6a2f3d0a1c72c608cd44ba2c257a8f2e06720d6dff272c9e180df38b460e51ae5f91c6339a1ab8b6a71584024d819a561a857059169feedfdbba2ecbde1eaad50c5b52aedb4e948c40ca2ed0;
    localparam LBP_47 = 10000'h9d3ea814195e877ea76de79f6b6c9c008670d5b13ec090ea284926e1b87aaf6f5fac35f4b2ff2b56e8478833846c014f4c3de80c80c88b262860617347a344f99e7edb71436f3c198ee35961b52eb7cbcf1dbabed302402cc326d6033c7ab4f2dfdaa7c8de34619cfd15b2ed3c09a3bf717e8dda40441980c607958ad1cb5e0d9504639cebeec5c77ea481b8e0c12201fb9405afa3212d0ad568fd3f4b340b531f015160768f0fa1bc615ebf4943ed9831935dcf97d70c920f30650e91e5eef0104b6e33db41dbc91cc7d553da7599770f142a7b74af3cd51e6cd20771cf208889cff59b56a36c65e6d0feaaf2e44840b69c714f54014c282e07b4e95cbdcf8684977bc6060f39a4671e809d228d2a669e2ed63bb6b87d27cb047ed0a6a841a983e0e1d15e4642fc749dddfe75edc7a1a0fa6f35d58261893cfe2f6a0b4596144528d0f699bd343d27d7ffd92199ab74011841ed06a0dc268269df0bf4eb50f3f839a29ef5fa49d095eda42678c154eda23b62d777ef23815be1f4b6047b9dac6f7e6de3cd9dc81581e331363954d0bbdfa033aec6094104a7cae847e224f77b470ff2779d683a1dc4b69e6442fc266bf4d05bef8b185d356a123a355524d88ecae61c14c9298e6555a16e461e23b35cbebf3c7951aa808ea53f7400c2b51f41c4856ab7738cecd31d70fafa19a0ffff12ea5293376fff11e546d23196b15f96e3682fd0cf81b22f6936bf6ade083abcba3876d5ba85934d7f660fe4bf20874db7b79c138007dc241be4beff97a33b3df6d84c968f298ab1e05144ee7f6ff44bae662183f09580e9ef0344b62042fbeb9a30deaec78e9a2dd37816e82be591ecb6b69bc264ac426c10ec9b2233d99b762d218fc14b47f8427d41a95c90811d2eab128f88381de5bd90bf7b99022682b6800b8d0ef9168fcbba1ff5ec29f506b375a40bb9148a5357616ca7cf41b214a604393157f941a7199ea783ec06118aa10952c8122b800d0bc77156a0d5855d0afef946fcce30f76ec2adcb66078d970d4ffc06e42fefd9ee3d5d189f14c4e85823a1bd692e9f1b8766d9b753356732af1cac60b21c9b0a612cc9f7c731466f3c881600b55b4c991d60105df15d0269de6f4461c49cb4da71677c9e1f6702981a1f7b51323ca975067c946efbd68be77b2f2a5e9a03f580d8c1a476f63a22f4e447dc099558b317dbf6e39554e4ef4d9275516c0fc52157306c8c1a164bc31d380bf4c28131083abca4aae4270eb3088a6619293437b5db66a1bd8dd3296ed0d950b31b678f737c2503c54eef30ca4d16c8424538150959d0652c409daa66b4021039227f24ae404226705d69f0e665fbae0865f21918b35d5283e75709c59b41ae6801c26125aa697db4a9854177b1290335af59a2c339ff6bde27d9743433c59f57aea5f2bd702b3fc0e38726731c22bfc912d83d152e79e13f32c210605b30b54196e9afe02978edb80fb46a15096c30d23b43527889ddb05ac745a5e5c9adf92ff2a59534214656738e0f31a5b74abe36b897cefe9ebc2f1fe2789d81122f48f1a6756d4e28e077f21e23f3ccb2f3baf31ab06e8920868acdf555ce65a3c1b30616d9bf4d5f203c0824fcf5004300ec3d071ce53224f874be9e7d698ec4cf683222ffa603432b48030172034f6e97e1b9d0984ae7ad6f71655c5117d23d1fb5f7b66469193b99e0fc5913864cb656a3cbb74e96196d7b22f74f12e67340fd3e01768e40a1daa8606f5960c20ff4ab984a;
    localparam LBP_48 = 10000'h8e27875ea28a8987886a78670623260ac7c577b1607ee62882ea3d70387543f00401c617053aee105f30d59597f3030a71eb286de958456d684f88d479d14c64edd67b1274a45beccfdbf3a256e6cf5c141d032939219ac9475bde55ac3366918e35a297d6d61f3bcc9b0df192d153b52d0b1778a68bfa2e0b773037a8a7af5c841553eb2f07b33c0f00729ddfe2536f60303e9e4279faa5fdd5a981411717dc3cb69b001a3a15e0145b7dabeae3f3b6aa6864e8e653d417230ce24f4a63afd6b5235ed406cb46cb4da2aaf5a42d79747cd64d42ee59124b0c58c717dc7021d4b4c895cfcd3125923529714ff8a9aad256dd8d4749278053c126bc9633ba691bb044e8ea609b4ce41c363db803f7b9f9bec620e392c1964d539f97340632a76e22dc9f245b0856c4e385b35a716f63605dc22b9aa7d9887fbe1621dc2747a5c3a1b4385be29334264e7a4210e59fbf039b84acd5102014655e237ad0bfb5525a8c09b6063a40fddeb8df62629dce88256f7c9de50e5e2c9e4e6181391e73323d6ad1147793ffe2f717bdced355235e89e776c48760291b53317094d471a512484c6e814a32ab98b99cfeced3a66e8fd436a95d6d8ebd6e68e72bb7791acdc0779470aefff8c1822752cc4d8b28863835e61cb9c7e218348ca69f13daaa3cb71e39ddafc7943b8028b8babcca9abb0013b720b4e68590ad8b47ebaa9c82252b637d814e9d37ce04a88a99c6052563d7f34f99f92266db7325a6e182ee2b589516650fc64646153a9e022f32fde88679247580476bfab20dfd1baa5037c83438bd8ca35210bd75147964a6bb5039e912f6ddc61e5923b8642caef68842250c8418a392140755936da77fe3e5ef002f927ba4f370df87e27e823808fc6677979711c80fc274c8818941e22ad28578b17fcb50ee3bd0b46c730ef12f45d47cd45c27922b7da415a9693fc0c37f3b2c7be6891719688e214ed37a1d8a9bb76c3aa7202abaf4dd831caa5b563bdf2166417a40ce50c4c671cf6f7d81ebca51b9512c0bced7588b5d57337ba4c0d8ac9c287327f2aca3961d2345a69a022682ee8f8804fc76065ce22b86875f450b863346b91d125c99bb94d56364cf9b672ed203cc74a77a0f2e31f350b814794bde43ad40d35ff2a25068f7724755dc29f3fb94c8f61ca83c1e9727c022a3dda76e9a613440b26b4ca04e7269c3ae91b24401ebb75bd5b8f28d94b8eab93695c698f3443de9f71fb804ecd8070e517742a8181e3e5352a97c9a91012c0b377fb6aa9298c804596009c2d2894a9452f740981c34df16a9123707a0d72002cc0ca8cbd2772d296487644a0ddf2464a9adfdceb87289f2114540c736f5bb2a376460182b0da9adb649069ca4376ecc1a15dbc6fad6af3a05b2d580a0f1e9b586afe0c7797b0fb8eb302cccdef771d05ef4f3545174af49fbdfae124b232bdf24d9d2eeaebfd79f444e768cab1c5165d5976bc20f7b94a8a66c704b8de26b7b38c2b91583ed2217c21a4c95f22eb777b8e22fb3ff4f6a96cd4e570cfb27885bfe13bf78a35d2de39d230611fb4e9d2be7c21b2a2638e788eb7a9f4c6516e99b0b737c5010cc6195b202912c9c47b9490a90301eebfc12c2a7bc9d3f9420abadcf1f1b993bd60f571aedc00c695b585db504e9c013da515eea99a8dffc7408d88f5d2110f2b291fb762a573d586ea1e611afcebc2ddc5139d893c94ea894b7949fdcdc5ecdd76aec3ab4edbb3d58d3cf1781b993c485622b9e5a;
    localparam LBP_49 = 10000'h292479c4f51d2834fc7cf7012e99d96e48f6e244e5987763ae3c272f296dccb9fa7cdfebe86d130a62ea380cbb1cc7169beb05e46b10c2ca31786a3c54767265863ae0391d63776308651ea82fa3145f6d7b531e407002307657bc14db33e84e0736c082a146823850527b3a0a666455e808e1622cfd8ff7660f585fc1055edf389619e3fa99281a58a7632a8cb258bbac16e9f2ecb95b64e57f4ca13593a654c0adf25e323f4d0eb176ee3bf17f9789376b77607d2fb616dd69402ad34e08de12bf35025979f7ac53543a93a7166a463a3ede11fe3310f7125c817ec8a0a672c50201054b99a7afe22f611bad036b991d6c0d0b79d693a04081a3f3f30c805c7969feaabaafae74b9fb4a7ee348eee5e7be48a782fea515affe5f9c27f732213456eaf63bc049c80d15a024343404e2b359f3985436ef3931d6afb4c5e3aa950e2c23dd642d8a4ba4e787960fe44f2daee0fa6062d6bb7c851ba66751436dcfdc786ee9a2c486f9bee131b3ce6d51bbb646dafd4626968f627be48b021b8572977b5ba78562b30e7b198dd013ebced66ebcb234dd412c60cb96c58eea1f9c73b64a14334de73656fce0e394c55556e0cc2ad490b953d6db0778cbb98c4e31c9f4de7c60c414a546d244330256364d116106297360cdcc7550739a133d0991d15c081c90b4daece5e2b31157f1fa8070eba0d39b870b8373bad4e51811d56454b226eb65ca2fdb5e6c75af7d445c28d67a51f80ad551395bad2b82cc6445c251de06299e1c6bcc230ee0c1aafe2527fbcc8976d332e83886292ca2cb62de17e1e7f2fbddf28018867501ae027cdf62e2a92808266c22ab1b139ce63109e7f64fd0d481e925993a6ac18e454b839300733b9af376d644c6e1b058b1e5662f9e6a9ecead9658b3c6e83c1cc25349dd693072e897d011a9ed111edfd5c50cc110c3acc9a77cd9a500f58712cf4d3558df45a8e8670fc93412276433d8d8716322bd8761367c810d1a697864e004fb462390249f0eafa708cafbfb91c18d1b3259ff43a81fa4d1871895c18ad0154e467e7dce430c8e593cb3a80163926f950f564935f87f4e95ca2646263ff5928ce5fda61f716247426b3fe284601249bf0e8189d9d3826e9fc47581ef2112cf4e9891e39d3562109d79b37ec578dfc6bbf5083ea63c4c4dc984e14103850ffb636957766642185f8b3d22f639f475f8ef8a51dbda3b968676d676d9abcd2196a661d783085dbcaf350bf1e94a1f84390fd770f11b1fb7eba9784313f78029ee6f2c88a9f646080e8f0375e787885df8b8e657f5bd43e1724b5d8081edab9e31f915cd44613952272dc9ab1c6a15be45625040c45f215084049e0e0764dca4898f1b1c3eb3e1df026cf7a8778d8935ec914f589c0a976b979ceac8d8560f7e87988c2d7315e9e61aee790e77c62ecdd7bc30a3da5dc9a2897cc797dcd3776633459c26ac58979e1727d50b60c6c453a24344881285723ce9c200537ab53c779e7d9d69c0498c35d918009b24d1e9fde86bda346b16fe775f89ebed7854ab34cb45a2c6d64358cdfa47186ea834d50a7d3b9073f4f51d629009d3741405dd049ff41a57c59b45be82574515511a68708328d9824f7e7dc81805b39d2d32cdfd618b1f4ad73c78934139f33a26b4b5a92a1f3217fbb49198b7b03db7a751956a112752c6de5f0fbc90a9d98db5156e0c9e3e41e23602568bcf7b1bda3985b9b36ba47793c9e86ef007dddddb5074ec2de32a4d16c3914d;
    localparam LBP_50 = 10000'h8ae4ea77c7a6e9715bd58a7480a3b6a7ccc80f34d2b7313caa96a15dedcf7b53244aef66cf64066b7d4b226e29e984530f4c680fb5126728a3b914ecd038bd8fd985f0ed30a69fc4ffe20f41dcd0b5567221f2bf67c3aba87370947602b62d9140d16ebbbf34497ecab76eaab2c22d9a5a42b907a8f41e4bbee04c0305e5cbcad386ac6b6c8604abe63059e44a0148622f3bffa0d33128b5f9144d206bca3168f80d90b36b5754ef5af147fcfe1d38a2ff15914ac70e76f33c37723cdf85e61409219461f3dd6e602df628be034e8d96a18eef1839416ceadb2dc37f1c9e21d761c63144663763b10de8a47fa4f084d6ff37a80301da01448674427b1f5d242ed17d19a0b61826f518ac52eea7344f232086fdcedaf528493ae2a472de9446d22b87805c5b4f0d869cdaf1d3ff320781506283809626b85f4aa75b633f0c9438fd4c3f22599947e506c0f78374ba4078189b415d4d0ec146574efbdd9586657dbe080ce21bc6a6bbba171ff0b005bf518b3d43bac87fb784448928ba5230e4f79d1abc6e9e5819e1d2670693069ea5b093f66d5510a3f7b8d4b429d9c60d590825be4869d6e231ee5074ba0bbc737275ad55e5f16b482e4e32c1402bae52b966a2e0127e18f534c373ef310c7b0d7d0251e8e397a5a9cdac9525fa41dddf51e9df04f1b45a2ac3ca86c1aeba288f1642d0d7c827fc689217f4b1a57c69ffc1cbd6a34d8e996f2081cb99f9cefa41adbb0b2179c18e3344b8145c88d339c7abd274724ef3821ec0d9e8a0c822722d84614a6fabecfbfca7dfff96922e95f9f589db0b7770287fa6765b660ed8b5950415b20733113d33025701107d46ad025cf42705cecce34a6a680840f77674eb9cf332c2f7c993a9b4eb8d199315706efb9447dcffa0fc452a1f67036b84ed4ac41b999ba98148c73da988de1a250e1c4bad2f7491825681c667f376a6906893c68c73cffe5e8b15a56a5d7f7a91bcf9402f29b6cc250a47df2a4c7ef80f59d2347072c20ae4425468dce0c16b49d809edcc91d4127b93e1608f88d4c8c4820a0b0cb7ce105e952f0288a4834281aa2d9d9f62232b05bb73372e295b026ee539f5e81e084fbf9a25e84511f48fd917aae87358ca64f9f9d94785ab66cd6cf4e3f3f3cc8920f203747f1a9d0ddb9bb0b9188e6708a959c5a547a70b60c339a19cd90a081930f745707d1da36f3d0a5bca978a585f1c32ef6f14609124ddf9af1cdee7f0193645a8b26d4986412491fbfdc18641c1086f36edd1ec283cc69fab747d73df2f30095d6543fa8f05cc3a8917b0349e3357a250f3d1c949152b76cd550c3aaf85aacdd0f2631f1f7c28935561d544777826d0d454426ac361a587ebc5c083e8c5da199fc881493ad276455ef982e0148f16e02a854b1d3bab3619b81f181d13887e30e2a451b1ffc5d4264bcddc3bb5f98d2de96ff0c3a784c004a99e7a6cb4b1f65df9f527ffe72ce4da6ebf56afb9703c5886bd0504728edae75f78fb7f62acfa2ed8441043d8e0786a46678fc619702b2f7bc161f7a7a0bb2864943c6a5080fe7bb51090631bf958880001ab9e49fff48b6ecd8074a9af6f45af4d841cbc8478a7c6c14e06ecefde22fca7db2c908afc20d9561c66c97e5fdbe91118a76ced82a5e9243ffafccf398605fc4176c31c78e68f8e485d34a6205df57e995ad3a661b45d1822e522f906ad57f57b9a71378ddcd640d46e6be7ad115af055c4a6eb64b83b44d40fa504f2cb763565662cad;
    localparam LBP_51 = 10000'h2c081089aae7bcea54b35cca086779a2a6c2b5debc1a73b8d3b870cd9f352e4df81a33ac44fa4f7b3330b69a215addc0b052d51ee9574178312ff2101209707f9c0a9d90c02fe9b9bda6a068021e1f3f9b8923ac3bb2808dd3d0a29a70e220714f871debdc63c565b4e1e00983badc54257174d0c91b75a705f8003b6bbea6791dfb9ffa4318237bd7e8f297439b231be812e14e6d4c8d81bf1de996497712f6c87415935cab25b110c0dbc97244d57553919856769e66fe7eec43a138e9f33a1911eb25f4db11b77f5c9cec0a2876629e0fe9ce3f5f195aa02be299d2392158bdf488aac9f7242669c60b464ecad8772f345491749be3009ad63455e24bd04368c5a4626f8b43093c2733ca3a9060abd6a6661aa2f52ad1e43d23f1b769414116f9a1f6aac1872172717b28e634ffe2b139ee1fea1d53ad42bc06452b87993a53536c45fa6cc59341d52f2e59a37a962a3cf9f8f45d4634f557e63fcd69cc255fb4bdcd83a6570f43e199d66fbd77f37d275050331aabe16e3c71b5a04c341ebe7b47f6ec53e359110253d7440267a79dc36afb3d0675ce2b012ff3898ba64027dfa702fb2bb81e7c1ae9c0373acc4e6e9d15ab5e75dea0a702468f884acce4abf6d8bc6ca5b4e039802fe9ecc097418a271572adf98034d0d4312cdd1453e0b57e4ce095545d48785400fdcacf466158a4c08c192eb45cb14ffabd8d9317650c6945a779011cd656c65dd2054d002dac9cb5fc4bc35f5d08cd575c9d59f927fef95eb945c54ac9504764dc8b8bb818eb910a4711fec89434efa7924c7eb647e1531129de849411e0d2914eb37facf145c1155b5f643da5d8eb7df4bbdc5b41a13a3d8ccb31814eed43fbece7eb656081d2ffc2277b67ede0ba3f9901104efc5d84182941a1fecb11687fad175195e82fbee978083c12af33852cb27db365628019e896772920b62ee9536211d3f1d1ba276a87e18a305b20c40f4cb40fb767423f6c154286d35c631d677f374a406097fe6d2fdc1f245ba334e6c6c897025268036f39db302c5e17640ec3eda9d009a8c48052385cd47ef62b849a2f79a709b0c78a150d7074806c37766c58126e8ad2515351a265c7a38e458d2e92ac4cd8e428466f2f46161dd912980560692b08501c37e1bdbd45d12639788962dae72999d0b29d60ac1117b21cd775962ef567b6d9a459a1f1b1b4247b5ec978bf72420af07ecf3faa31763d7d741c9b17f2ed7bf490da12cd59386d235bf7ab5d10ac8db4ccd87d5c96cee67a5ca19dc61cc178aeea0be201312a31fc67e23b4c0cd7cce1707509046eb382d72f8c8794ce7ae951d940f257b572f752ea6125811be7dcdcbccd376f0f7136f33bf3065289b5e137fdcf8a64a975f25c8465c77cccbafa6addc39eb3e002af2c6d112bad89086261c98d20f7a2d6d5149b0c7c12cb2d658c91cd258fab5893d3a80825470e6fb5853b4b9ff0d97625128aee6dd7ffad0f567b9e6434d931089e35d8a012c8196f3efcf901bbc8ea34bf55451d7834873db8d502d1f44e5ece6ea79bd0d5dd596554c47a5a6093b51340f39bc6b20f019793adaa70b12b35877b3372e328a2f068739ab1918b2093ce2d2561aea4da991ff03e6d5dea3f7a040ac6748dab8e005f55bf4c0e68867156122849e5c815ab73615a75ff3d9a93e6a227f4d5e5ded739f70cc41676281c4402759c9380a3a862913226e405c3e9555f5e09c20f04ac974f259553648dda8522a30b57b7dbb6772a;
    localparam LBP_52 = 10000'h7ebf064121f43d6f819ea36b6dd5c75f8f96e3680a72714339ab2072e23af3189ac8c07ee8ab526afbe33da565ce21cff29a27101ba98e6a5417276c575546e1dda2822b17ed624d258a37c234829a44ac1fb015a9703018d80d6ac14e4fa0e027e936285e2614a0c7985010bc34d3f8f091d4fa6d0e371408f1751541c7d8fe8393a38b4a77b8e4512d4fddac2018a8c3a797662c3cd0f9cc148dd5c1361954524f7df24ee0ac28cf5a4efaca9783c762abafe109a5ce7879c7e22654d97ceb30626bb3f3b6ce4f3fd0a9d6be2688ddc17d17bb6f325f4e093969f7c7db78ed25bdf696919d62dfe321d6f679692c4bbd22ee961b33b706dff611dd033e86043889cc9a223f0eb4248515ea5b25198990da73f7efa41213984a0c12a0179f82b6e0cbcdd2a5d558432bc1ec94723d8b17d9111b71fe583bd1bce74a053f831488ec309510502df18a82176f7589d4c0c8fbd57baa642e8e79b77dd99660d4edce3b21be3ec8e271463ef328b648a06943cba49fc6b56bcfb92530e4daccf0000f862d5c4a23e7678035a690a4298e73f80d7362aa81041d13748dedeff6e5fd8ce2562169a991305dbab68f1bf7749d95534b0a7e283b7084279f1156844aed16c79354e6fef5aedcb158399c85212f2fff9b39f7d7c82d7eca9c3e019318d11610936e8fdc431bb9677d2ba11ad0fa92926a698659476b4b8625b575f845c3b4260c8a87be59b8675638de2c96cd5b639ce163cc1cd44271277876cb292734c2f3147855834a44c14758e9bb98bd7c9950c712f8acd9cc4b7e4c6d87686c66a1c611233bed046d92b3c36f5f62d9306864abb4c052d21ffdc2edde1025c13be5c00b4e54fb95a7bc0d23d92903ce8d37710974ddcc2ad686f37e1e921b3149b84773d62d35ccb7c98985bb6b95374a653bdfbed0c1bb5ff865a2ed93142f7c34662502aee788949ab3042d904a79092681fe66a5bb72c2b2d5289deeb7c7bf66618bd1a776e28488e135d8de7427b8317defe0228f94c157e309bcb42d9962bb2214120b6b9e9fd856ec8fd8ee6a07e6cef1f7344add060d5b3981594a7e933f4e951405795fa919fe6f9181d1cb2af931cf5c262f039e43dd345dc34b19bfe0d77c89c30240fc5f2848cda7486bd5302add9a478069e60d3527674e905d6b23e39a2e4dc69479aa36e44b6c79c375960197de9a63f1dd7e3914bcc4b4fbf856df69713ed41066cd22cdf27b9ff30b0840717bcffdde3cde94c5f65df094a6d5080e10b38a3ba2927426cb52cb3948efcfba9309c84e3516a62edeb0fe8226c219a3d9a339a0aa68de58473562752018aa03ec2a0ad5a510c82673592b02284b060656bad16004503389a1dc66f6630a649c73c1a7ea53bf0d7427428fd66987c1342d08229887888aa6442d6ec14014bbf545bb07a44d982141d4f606b714167fb3352303c9d621bbadf2ed82b0fc1706c3a8ff80c7494fe561a07d269a9f370713b828a02979c4a086a7f5dbf2bf6507942a1fd481a06aefa08462a1a50fb6319c435f18c9d3f776a7cc0073c81ed4fa56f175f4e7ec17a15d3f290eaa4ef1a694a534a1d59a3d803dfc3ac62ef6b265535c64f2277cf9aeec369ef3ddf8c48377ee6c263bcb641dfa04d7165e84081cd130f6034aac3395e41c26bb67770b52b912dd1a094cc40b6e13e6cc35cfd156db43a9986cba799f7693fd65eb296886e0531b4f5dddc7aaf794d06c104682ebb48ac9e95410a55a721741d52a383f39;
    localparam LBP_53 = 10000'hd7b070208be98a35899802f63ab86e82ba35cf557d86d31cafaacd4c570bf312a77663c48b1ad862cf0e6e59d45ac7328d270104ebe92c567bdd05665304d4cd4b7e11bdd7c5cd29207837a2bf4d1b274b2ab277b43237476db51fe5a690e78451830d957f5cac6d25136836e194994a3dbcb1a1fe7b56a810b444b2351a580e1aaf67bfbac96ff506f69e224a714c5b5132835e6ac0bc3a3bc8fd4c8fb5375aeb8c704994ef23a6dac2db43389585d705e0d98394268ad13c73223c1246adb29a6d08722a1bc9c0ad2321b47d67a8383d72302dbc04db1b36d1d7404f6ec459e1cbad56662718c683ee75ce758e01cf04b3744554b29c55bb8de0c210928c3642812f75795e6b77d8793b3eac39df1f6d3561110ce0cff1c8858ece8165c22e53d0290fa36894a0db87988eb4cee405498a0f4fb91ae25e736680f20cef64021530ae7f595ae22dc026c778898fbbe64a8de3557b4a50189904e1075e7075ecc059ad5e00c4aaabccc19837712c25f254070de0b9703c03e36cfc13cdef3dba844b055501cde26be26b8abf4e86f8becbe22d1b23e9d4fc4541e10d5292279e927c3bf38033d4c9d87c481bcfa8e73262a5b29893c40a944e5d61b95970e9291894d94e88691c478a04cb996866ee9a098f1cc374b89a26db419f879cc3a355711d7ad63f3437ac8ca18877cd5b0e71c29c14338712e895641b698b2962d6b8c63628e650c7edf8c83eff6d3c531fc6a5a6ed95fc7f1d1a343f36fe41d476afab3329e0d04f93e3106d03ea1a33bda5a0f44ccdac26b5911ec8f0a75e9ab80dc8d63f3fc0ae366fe5a71b30037843f19797dadfcc636bf371988eb6fd2ab5b9fb18261c4dbcd2a68a1ff9231c63a0d3d5b136a4a85e1ca10ae57764e313bf85497a6e46bfd613ecc8066ebc08af90b5a54d7aca2868e4c2cfe77510ca212a7dff0bfee9ce9c4952990c0e57708c8855302d2e2687d09a83c20a1126212311bcdeb44b3a4e56fd6d546a339c2fe1737885f801bade5788ade0580db14b770dae1c14d17c76fdfc95453f4cc3ea11e4daed16a8ad88712ee3070e5039dec7ed6d08061322e08d9262d527069b99376ab129c6b394521822c8ac6193506a588c7643a1d8177d12766f34f40ec135e8c668889933760d3ec2cfd65e24618df1ed0cbd7330ac219daf470e954dee74c6745bd6dead5f71b7531b5ad438042f370fb54bb61e51060c4d0dfee7691f3f623ee4ab1a075accea5960a7bbc1cbb39a4b84b840c37879d6be1ff1e175cd94a586151bf83653c5a26a9116e9db6e712f0e8b97238bce1f958f6d365de47cf3ffec70065fddc13620624cb50fe8a9eaff27944495546453baa0e146a5ff30a96dcd6b2d3ddbf57f2a490cea2b22ad684fe4e491dce340ed7253523db8299a08c4f52c1e16c1afb7e337aebe47fc32abbecea362161cbf85bfbf830d883b0463e29ae3d3874607258732619ed0a98ac30d4212951966b1ee6ceeadca28e6967f3dbb4a1e66046cd2ee0b252dba147b13a9fb132e1191c864a55f3116b4a3c1f550016016d3ba35c3c3bae83bbd143f707f2d071133ab1e5f9677c4055c653a5db5ed133c31c47d1fb60e3368fc8e349c6eff0fdf2c7b09f95478141cb70c4ae3668801e943633caafa32453b8a8642c7543bc6a10132041d67466b5030f9e8ac9fab63e2974c54bfabbb7e8b9be9f807f9674ab5b0da7c7ca46b81d13bb0cc7b182fd85fb35dd6f441e96ee452843cd71c024cacde;
    localparam LBP_54 = 10000'h748bb91c4b7fa4435113c5ed656441db3b4e9940dfb0bf8bb3dede991ed1058a1e33dcf1315c7c19c6c635721a6864f45fb11f7790b23ee680c1d32f171bd17012879d1f854d44c1e646ba3cfaf27d2a6c1cab077a686b0b32b6854e32f5c132ca6dda77bde69f12a0678d24cb055eb75ad5a703c2aa087b42f6940f6a09b1fa71f7b63d43069ca3c22f47b9c051b77dcaf33adc07c1f96050f738df05fd72a6641c588f41d782aeea4e776473d1e55d4fe7ec9bc79f6dc10ad51d6c7224c67ea386946286eae266e0883670c2dc188f8ebf4727adaa164567540b53eae7209461edcca60d22f17dae88a104cfa02f0c7fad5e88f89ad470a05a952409e6554962acf9e0f4141ef2e77da7847faa8c2cd71921181341be29ea0e27566189671ff6b73340910c9544ae3651d6756a654bb9bddc58126d8edb3f8c0c319278c1a7faf35d7a5da82da130143c33295e622998db5448293d9cfa6e03749ea2f5970722620eeff9d349a36edff720b14d025901b092da9130b92589a3715871b74c4ceac3eef116b39907f6a03fc74644e9f5dc3cae7e13a9cfb95bd396bd6f3c38696d736bfadfb0388fa96395b64a2b41082705550ecd77b1247eaa41c2b496a5aea53a0a6fbdba108aae932d51aac48cf3e0ee30efca12df2b5a34689eca7f0bef27477cd198f9a139dcb66a8471c8e490af1ed471c2c5251318455ac3e993246c779d9dc5179fc5a3c05806b4d2f8441b8d9d5ec39c8aee05240d06db0e2992759981798e2207a92bb5f40cbe53a8b2c1831b34bde6aafa89bca9c940803ee07de0f10f2db24e0231684ac0918f7abbf7a635f6ace85eb9b0935969a5f324954dcc4b87b936cec72c1819d479902afce9db1db1d24f4f63f4a5733e0f238e917a0660ae4ad62eb4e03078030783adc6ad435d8331890275099e4ac059330b560c2cc88b69ba00f3e062bfc6a60bc3bd405b766562d16e2b9cc253576a3b6688fd23eaec3dd2631377a535322cf73bc9922e92775b73767f7d977305479c5a1c6a4718ae2bb5d9b4fa1c71ebca9ca2d9df60fc0b6644afef80a2e119f2f622ac86efe32e0270338dd6fb156c06f4f42ac776e1c5e0a5a6a1d90a045d13dc686559f76955e521512baf1d54037e1907b3d19527034eb72ca0b6939ee51fd294daa0598d8b84550d568383911ae93d48701c4db35af27eb56489d17e731723909ef1508a6d7d241a9799165c14e8416c34a82f442aad4899fafec36e42983d78d6ddea34334b8e01fc4a1c4b41e34500de3d44fba27491fc293564ccfbf74a2db4269458582dfcacdd6a634e63aef372b1e8da08ed9c779893218dff651bd30fc46b8cc378b437ea70808c12faf86ba823cdf3a8c92c339299f95411a7af6b71eaeaf7302873144cf958839879c0fe093a253a9e69c820aeedc893604032e0ef509b6ee14a80c843f75e1f851093d50bb1b65cdaf4001f8d9a5cbe21570f543288be48580a66fd41d14ba5fac9aa1842d8c2470d62eef25a707b30056e70ffa53979b2992d4ef291212a2b36ff8f6baa43ad549f1ff1794f302006631a51fb9673d6ce921ea0d326638c1e6fb0fa37ac8d733274be95c689fc553f7750225c35812fccd8b29d1ac7d93dcc831781193701df2c381f9dc051f1a9cd9aa5184523f1e56ab476cf5cc349107b74a560d2cc42be1e1616fea2f76ae840f8002b8b36775d94fd16f3914ee30a7d4fd8ed50e79d584cc5ffdf167af863b64c42305a8f7f0b84dd;
    localparam LBP_55 = 10000'h155150f68b2c03db2b667781b245250d4c62565f6b4842ee92375272714d9f74cbea213ccd651291a1ca6e17782418ca7605d14beb4953c8394090f6b39296237939e4328cc4b12fc02841c40a024543fa61ba1f9a999f6f8b9465ba2121ecb302c7e0d45705eff458edcdec8231dfec66c195843314508a20c5c28da7ac67ada616bd3e6f704eade005e324fd970a2406dbf25ddc4a5adac29b75454183a0f969c4d8793f3273422b820cb51ed55e45423b46dbc186f5fd801f14704cef357d324866d49030c18b64f91f820954aae1c94615edcfb28ff3430c6d0d4e67797d649f8b5f9adc630e17a07e9a69591f31bb02de598e1550fb14a2b918e1c56386be7ac4db2f6f4dcc3ca0a76a1f848ef195f89571e69d70204b5e60a6e1f67bdd9b7556fa387157d8c0d072ca1c1b7a84d25335554f73366dda7f62670e7ea1fc85334f97cde5272ada6d3b9cbd274a079b6cbcdf86fb07c0db849ae73d26fecd73a92cbe802331b1dc5bbbe0ad3519ee6770d4fec1cddfe48c4636e6383666b99e26b5072f728b03862aa816ea3a790c74c2489c6cdacb214d6d4c1941cd5c2540cde1dc3c61152006115991562a8be7da64d82b596198c1c09c713688178234271069836ff265a9d3d93250ba50dd96ddec12e80c14da715231f114d38fc42ce3c16318c7fa75a1163aed46aec268b2ae55778b938c6c8f515a123700913e0c24c20aa093ce4906c9cce410b5ed82a5d181aef31d9c56243f614414bce54f6a4ebe06fe0be98a9fb31c389153779928f73cf13032ebe5f903a8bc88bc9c9aedb6b63012c0a11c0ba86b806d36c7d3db63fbf55ccd3d6cd79eaf4b5475ce1fa02fcbc9c7c05394bc6d0095b21d2ef5df326c976eda4534df0d732572959e80019ab59261eaa6754832447274fd2cf65c455f7ac2dd7f4ccec18536b215bab683ef3c9a78232833a9cf1591e2eb569de979b320dcc29b08b44caadad737bd4dbff7b358a2a42b6eb5d7616636c70153d69e6ba8cb9a0e90536a6455db60bc493820d89afc9d45b6318eb521036ba5bf92de5b8687f03ca58615069284e1cf8e5873fd81c52dccf349da9aeaac1638c9c441493be6b4cffc3682fbecada68d36cf1b7ce9bf64857bdd11adebb5169916b9c0082c556a1354d5dd71849dba80ada5aa82354d7af8ec38118f77bb9a10cc87be46e06100b89ec25eea16c9327476c0cbfd3c50a57486f23a64a5dc9bf3348dbb50fa12e032f159614b29059409759a83e0ebb3166e0bb9b9c1e79701e759378031b96783d024cee66529871eed2b91c55ba4be44fe6283f8dc444dab6ece2691f763ca45deae4f8961e0a84f5f224535a5f20c35186673f38c29abb07d25db799a7d6c374b38364f13cfd0deeddb2679a2f511e31550b4b506de448c3d9f581febf44c49b54d8989ff0d0fdf930c29858a378dc73e6c0ce991e21a459588fd261fc69b2d91a75c3083fd2153ee61bff3e359ed322fc34f564b7e6f51bb98ac6b53bd2a0ae64f992943e20d3339681d498a1dd3aa0accb24b2aa47f243b8f477dff78499e9686e4ad8b16b2a13123cdf72224fa1ad688bb759a3f556bcdc8269ae854764a21c0367c29b5abcb817767fc947c28867796f372310a258d1e2273fa78c14e05283b191a9bc9687abbaa543b0559994244299f3dacb6d1c032d4378d13e32fe358f3314819827e76c095689e3be5f4631583e7e1d58ef0b1ac36c9f5faa8ec0fb1fb4f59106f73d7044530c8fc;
    localparam LBP_56 = 10000'hf3da19217515b1bea24c97f1fdc58f067d4f38c9a65cb5ced3b767902d9c90cdb9b012a295706a33b2df965dd99ead6dc5dd5c1a1a7aa098d1e570bdef9f210fe40d833177d52c1eac26638818141cfeb23b61cbe4bbbb685a524134ee17c785ded5eda2a0e8a6080c391b3f499fd67c1925bef038e30ff4abccdb0dfdfd1541025d089804f909f32039564d359b381aff0f8aa55d963dca61f66f87721944def3249ff604a6f945b29c037c74cd538c709b6dda5fbdccd127bd18ac2909298837148b1bef133f7ddf203354cc7ebacc3bcfe2045c0417c26bdb0cdf698dbc72bc5d47e96150f5c9e64c60ce28870d601d8a5872093ea1f7d4e4ccbf300e7abee70e776724b5ec2c94d248335f2c4db08b468c1045a44feabf9808ba314db7b6c697a4b19bbdd289cb169c63aac07172442d2d651efedf6ee1c18ad7dc1d25a0631a1c30f82a122a460e241e00b28aa043a5b1544908a21f4b8752991e98e41a42c14bd356650514d9c85e30d86d76f848f68f90fc7dac1579c012679b6e76fb838aa6fd785947d31d772783192710c8a73258b7356d9f05c85451df217c687131b491c7b76558c9eb42ec47edff5e56e61c51435d34dbf483fcfcd2d4d2f83a4459367c257292f400abf59c1fdbd91b2aaffb148e16ba68c1f429e97169d1f719b15b93b5b00b010f282c76ce8d61b3b4a553dca8b41f2a00210e0f7db2ac15167fe54b71227f9e0707737877034fc3c52d24238965e1ece96b281134c3e5e0ce6743736d05536508544816c258d53b5b589e48b00b2197967ac96d97d2c89730931d0a7f960aa8eea430ac6d30f79b67a551a9320cb2a04264ecc42aed1c1942817c3bbb4d75ec2a66b7d052e6413f6537648414652fd0f7c533d2752d6676c81983f08e4485ae1c6b1dedad718b3a749ea9ea7a0f2c30396048cff3df10b60f9473f2b725fcb4af3c648fbdb27891f334eb65ca8de76dd102ce0db8ab2a44bbc276adc6080b74346dc42bd2413f74c2ee42b60e03622427407d96804a008091f295d6241e9ab5a18ede9d448e624c3ba073a477d9104bfef3527e850d3a0645d187e81e2b32e62914d75ae7755fd072c0678e4f50ecc80f14cf1ece83345d4afaaff08be01ff9ff63923d85aa2b7bde2a709e07d5aeaa6d5ad809e58ce36af491173ae0adb6332fd3abb170f9d517639b670abcf5b90ed944adf76f266e8145a1c287578cc520fa21c05f7ec3786116bd276a87c4e5d88d0520f25d5e0aab60c64ca5803350bd6d766ff0645042d2ac2dad9f68055bc516194f4dc597cd4ef9e651a2da23f09ff93f4d27796a3e6dbc7740d8e6f629f7e58e5373367ff5eb490bda2cfa12d356af067d97833ac7d956094b2f8dd605eb79d3ca580de9ca85f5a606c8634325e071527cebc697fea9e20776c4c834e95e477acb7aa011dc7da280c0337cdd4b6d676ef6b7bdfc6b2ed19d38ea10b440561419cfaa0e00a26d097952a789fa880fc1c635de9c23f0f40a83cf6c69971aaf738afb90505071b38e718b8e4424b839c57128c103ef891f0dde121b5ce20d7575d50334729ca5272915b9a3fd5fc1aef28a8d4c694917a57e1400ab75e34cfc4905c254b31ee9052255d93bb9cad173a9f96f77e1c027f266b0e9a33547b985a9e21de3e9a8655e1741821b7eaf90f8bb956e63e3521e6bd7d2cd27a06e20a2cb4956ca47d62785cd81825cac710f3ac88218b86cee6fec73812e14920ceda958eea560492e7018637d;
    localparam LBP_57 = 10000'hac967876454e26903f09478ed2fc48265db61928b8e301d5bd12639052c17f0668604b058c795741750bf65b7a0eb635ef169117c9b2e0f9e3c70a96cf4ec538e8446ebdd43bdcbc4ad949160cfd5178d91a4ddeda0b56c372df7dffa874b068004ff0562afb29a55375e134b528d28b3d02caa84a0a892324af7a0772c8a9a0a0ec249d6d7a0ae34a6d26f67145b2cd3c0bb23eb7725ae315574ab7fb8d301cef277833708b871de6144579c50c4d3fc8dadc725acadd78bec62058d58fe642849f0796f97158c16dd79c82b64de6909a33dc938adc7db55df3e1829f213d5a5a24eba61b085b4bdda20e5ea076a6e82727d97c01cc4fb404c31a64e247642688df51fb4841646b5275b1706c4fd490191d9735e49aa9dcfe518b30eadb1c319db0335c64a2ec1f483701796bed65284a0ab557483120405d9537ae34f04f9e9ed679a76a6d69943f46fb6ded0fce2c44e3f00e1fc4e954c3ec52ece9e6985cc837bffdda7919351251308c55ad6cf73bd725cb651fb118c9e88a76d3e5f207d0605381414b5ad0acb718322f2a7649cdd0d16b3dd24826e35f06c8fe665a3f0d30230c04b92aacc212b6f0e895c5e3f72a276c3585d1f9ff5024e83b53aac22266ba07569a468025cbbc58445afdfda142d1b5b89b321176d5a7d487e6338d5f511e8844ac4fdbdd9470a25a25543611a978cee3e8144bb8cc1ff93fe038701c0672e19b9e4dd9c17efab0bc0b488bd1d8786dec8676d0ef1f1bc9571acaa407b85eedab5f2a7762a7e369b50776d7bbea4177eb08f624bba14fd4a6ba82bc80fec3901d7fe128a47bbe5ff656e147a0588752be1efb7ead3b2bff2215045c45b7d6178ee7dd066597b9a3aa4b11454d7f1a9fc0c0514366b17295e8e2998874fcd43ca51f31027ead381e91a1f38368276ed019cc36835bf912e5f8e9dd0780490475d357d41e80552c8f1e1c685d0041aa2c48c469ca99e01cfd43d65cc49a0ea24c67f3226f7e9845626699503494764c03e4ad5be0e8388635739a46362d8e86964e26368a8fedbebb5c9d29356155fa765e239e4abd7111c2456f6f8b5f445777200796ddbbd33149c0b09d74dc641805cd839f45fbca3b60c40f404c15683d713391dd83d79cdbfefc1897ce3550dbe0a1fc39f9d421507ce9d95d695b713dd84a38be1f7353b8736970514eca9e94cf7e3802cd67eaf08d850a16abe38d27327ee08eb98ce2eebfaaf8fb546eb5ee5dcf6484ebdcfc9bac45b2a63336f3055852c839d8f3c9c450041b4ca845bb0a4311a920cbcca04c31f329ab3a1e6f0da7d492c807bc264d86a9a6afa499ac4e2d4162ab55030461595aeee8db5b87a05b875263dc3e182f7c78fd08694103d56309534f9d88e1743ccf96ed849361de5770311dc0664e6417b79098251985aa5fe0440b3ac67676f05ea281b728bfc71d43a7a8f16f7bf01aa94f49f6250280eac2283e71c5fd8fbc8ee7ddb166a1ec50f93c47652d0b3b5b4ae220a3d9367e09770a78466087b57d0f55edb7262afb6bcfffd238bb2498df2c69d9c6564175ee2ebb37cdf6c89da07d9d86207c8227ec96f1187256d7f037b5d6b146991200065c0c30766696af1d2801206cd6c8d0511f8fb92eed85a72d10303b5f4bc08525520e83b3b18b1a8c31fc5264f2a1bae473ac387304ed90eaf168e0c560ce0e7f908db50eba86d80b2d7ab45603c60eb0df57073097eca6d6f405ec75497313afc85accdeff1ddbf66993f5172a38;
    localparam LBP_58 = 10000'h65fc8f434909bf1a37a6b0ff6a5f1f3449b96415a9d98ae8c9ff3b5a839a15f182a8154cb3607fb2c575285a80987292909a24aa9699bc8b3844bacf4fdd560a72a3d566591e28f0b56d45dc389f46cc39508b3379394ca3f4e8abc0bba1dbaeb6d240b914421b77ec43ee8a8aa8fda0eae196eeeb5e05cd9c331c52ea119a2b48861e43f26f5f47549a2df5967c9f1a05fb9cec94134e9bfc687d04d7e0bf6cd78fa36ec77fc41597f4cda95ae93733ed1910ba7c3af8785902c449dac9c2bfe0470b6d368c6a906db877798ebce44bfb836069861ca3804d04e74f3e9f4f21bf7a42ce0a1892f846061061dff548f6952bb2d4453bb0dbcfa10acb36bd94ccf9cbcec251c664ea87acd1d9c28d520c2552c84a42d2a0f8ddd238390e1626b9022c2f98fe39ca4b5e1f2994f4bb06db2b162bf4c066cd1c06cef0027c6408b790ebe22f9c3294e48cf55f53e096ac527fe7cd65000e21667c54206bc66e1a5ba78438582b379fb399dceceb58ba1ce41882779af4e31bad3887fddd89a275e901f3d0ec7dbbbfb17605f32a0d606c3627bfa355c2063e641293cb8d5f2a47bd2637497673f5ba21243075daa284eb200735365529395ccc1747404dbe803e2dab4d178425f635fcb39b8fa10fe40e97b2a5c77651f26cb31e867c313ac56de0032be3476159ddb5b965a6854e983965775d3adc46da04edc02128b2720a2c3c0e05029ee897bd6d7862af1e590c98161fc1546c35a614a3557edef931d769580c1ae6e35534b7ccdc91f13d0ccf99a14fffe9650caa021460afcb04571031cab5ecb02e281a59571c0a1c9aefca2daea4db080712571dae71b534c03a56919006b7366709aa3f811ee27e255e21f7d804e22568bd106815d2d5c2f2eaca76ce942c3e6435fb596a08c9bcb0c03bf2ca02d3fa71bd3b8210354da7a702bd03c06ba7fd6fe2c4d1102a3ee559854e72ee251bd10d4622e93301397c8e9025b12a1edcbe1f329e36a2be35c4270267bb4674cc5c75bcd7fca6cf2f0e3f5ca36620b0b2fe9c22a66e1a2656a1d57feecef20e9f824ff70e733db28e18a6bac356a9e5f582e08ac606ff8c012f485d1152459ccd981fc6d350cf89c8e8b683f70c2b2b75bef56cdbea8d0b113dad632db67204b5be419c6b7092991792ae3b7c197461ad8762fe14fd64011d8b0e777fe936bc336c81065ed4f337e8f930cbb6db8203b46d1c0e571ecb6ac2643bbd01c12e7ee4312101b386ce0e11f1af92227d38e61d3d67b1206b6f87c2121f88914db9994c74b775ef1adcc78bf3ab3f8e9a738831d0807d8d65c9dd0a180b4755661f59e78141f051badc2db8e2423f7f1feaf2dddeb58299910fa6dd80a678805d0419a50e06aad6931f3a9aff763567a388f6ec7b013c60326c44a5340127922473e661882cc0c66c144793fb73b7fc16b5359be6afc349dbedd6608dd77bc211eac2f3dc28cf5995b1ec57fbfd4912fa13c500ca32a102a77a58d4708b8829dfe84c5b14de61766e116eecdec5829412a27304a0ef33c11b141107d279d1ec6db3ad7b0037b404ba11e515da231428e8cf187482436bb5dd5e466722551bde522f59410100daa90027f8afc49ef641c036ed1dffb3c0e1f1a90897ddf789f4fbb88cbce7619c6d62b7c1deee512c06569cb6e217f7890a994b60bb6607836a06bc1923cee6458a0bbf85f56f63a462b05c3db7eeb34641f738470a4fabf3f51615fe1b5386c560782fcd74387b2dbe942d9ea9;
    localparam LBP_59 = 10000'h1eccf2da2102cc5e319cbeb4623c49e40f156cf655521d8477c85de066974a8853d95cb412885b0c95fe6dcb3adc4a52cfb030cc1bbb5d2ccfcce283ce5388f2b08e321abba5a3b6c2ebb7095647bc281e04ef9413674b4cd7dcb4d6b705d837f9b1d292c48e735db346b5b78c8e975951cd88b88034062c155c5a338e892f569caeaa5719550b270b0bfc6175047246c5b6c865728582f5c1afec5da7020c77267755dfc01e4cd522acfa97bc8023f9f5855888b63d0d08e6083f063965d28032210ec5053bcfdf601fd3d74fd6bfa55d5d6f46a6a6058fed02530f3d7dc96d885ac99cd3dabafe8958770b65fabe50570499722d8dfa7207499b51e5dee7d6e9b912f9dee6752f76821f4e3baabeaee674289c48ac0ef0d045123ed1f63bde14457bac00e3ec31163b31d724582370260815bd6a8ec31e1130f02341359b90e40946327b93224e17fc6f74ec9cd1b5225a6390160604b43eda349ca21858733d91f87184fce54dad7f1a0c3bcd9615984f3cc7a3dc85804cfc1dab5c3ce2a0a592a141902e3f5233e4a66094e41a5429a9a6fb8cbf14d0072f48acf1121f8c278bddf12ef275d731cea33cc8b5a5c12b688df038373843d70b7290b353e65b009b9f70d3d4cf4eaeedcd3643d1b888dd0811ddae7034dcc5d0292e5a59ff40880719a3c3e5d7d4b09e1085bc7e975aae02b03deaa067f165fbaf7bd101f141e4bca4ebcb554161a4e95f0a111815c6d8758f614a3cdb949b7411b87ca7c3f053bb1f3fe7d9ba43a019f71e16534a83b70c2cc5424aa2e32c3ee58deb7a730c0ecda57313a270d8d9763000025cc73b24fdd01668ffc55c3c7043c3813b4a30d66b27d3521f4e08f8b57e0e8a865d691d6e1f3ac0771c0e37b79d616321d73f81a119b6e1cd0098ac17d390367a1855f03d3d24462cd5b2882915bbe3e12de5a93557f0a8ba6fcf72a65701f524171163562d10104ae8a53de6ec2f6687d2166726bdb912b90feebd248cd4fd9e49d1b5a0cc64f5d9973b8592b070ae4034d4148d5e4cfd7140f7aa8947cdf054fa66438e24bde8d926196a2129df4528d71bc000763558b6e93f2fe9ba9953c890e4d47e17edcff4a190cdd442a9d04014559a0f2bbb77462ba3616d4c33eaf3d85a25742bb366baaaf3755a3bc704b1f0c2e50ddfcbcae4585ecb691ceec60de2a2497d5d07d2b1ffa20affcb979d39871117dd050bf8db8be899abee83ab1ee9a9def96b73c43ebb05d798f246a00dafbf030735eaaeff25a74d07ab7406dba4776a1a54e05a72eb36fdb1c38b652639e4a122a7bb470e3c3b6b91dbf73eb0e49bcbd06e848029aad328484f29c6cf1f55fb7817e7384635462e5d6ca1e0985e3da120340d182396a43a2036ba0491a3b6f621d79687fe989d1b198ec6ab7a864a70c59cc50afd73d3ee9a64045b4421da55ea7dfe1b83ab1c501068afd6e31b9653f77ffc1f6867e4c9d5e63be5c9a97d7e3e1d21942373b7516c6fc48a7a22d258ee1a9152994e8cccc180349e731c542f03c5bba2e2371aa37a98417b3b4c0e975656239aa305efa8ae98183cd59ecac5c2c689e3b13f6e5ae6c351101f5af27933a440aeee37466c4c7fbb2a841e1d0ffdd4d5a5dfec370f5f0f58d64d4a185688429a690272baea9fda1805a478fefc21d01099a3f8094f03152073d0c7affca12776e12e241f57ee11f37b8b2778824f85eb17ecc5c798346ac875a1efc745c54f4d1e30d42505f0907c92ab7289725f;
    localparam LBP_60 = 10000'h4b4c488a7306b4e68b65f156d32dd7a28f7a46b22bbd5b32c72cf06e75d2abf2605781ac6563d1b13e665d39840d3df2cb603938dc9e4a3f3d3c3fa371f949b96fd0c883e61d7cbb866e6f1b1f17f0d5b5fe24becf3353c67cec62e3afa95db0cf1af7c163df9aad2a39affa1e92fd53330a3ba2014b5d69825becf911ee4bda62e5f5a669ac39f755b25ef584bb2c2cf1f4af3459a58ef3b6d547d7638d6c433647d035d3fcb3ae221db5a579c18f083051428f4981e97a71397b4f7a8a3274c68a5021916390738bf92640fa36f2dd0ebb5dc3a6ef62aae3e926654a099c14d7fb4055273adb61a8655be3cd1c3185a41539451fc91ee0764fd1984035b2ca60fd9c8cfd9f6da0814c148fb5e93a6b3a062c46f30f67a9ea3dd90ab07c121790626d83fcf546dd0093157632d9f61627e1250a4ce89e7fd6d353aabb12bc1f48ac96e534b1e34776482b0964a3f05b98129a3998b4dece507830a745464315b87dc278db7b767ce7537cdab6e510ee52a47241d74a62be5f68452584759856a5454da37f87d8aa2c8fb1cefa1dd183f8ba3cf6ac39f94cc7472623bdb343a5ac08700fbc7df282ccccd4d87cdc83cb034ff6b70c5a0c04245d3b7a36d35dd1c4c87c83d8bfd4f63e12cadd6428b114637913f3f0df14d44a4c34553c2e11f5d6f23a0a9b7747a414217abf5d81a601dff23e18941641f829b7408e424be5ca5e2cf57000defec7976cb47f65ad613070615c8dc2a15211c244738a53eb9fea4b807a83115dc79b7797467989382df5012349208e78d834785a421281210e33f8c441676f5804b95dde3eae66250bf40c8817713f92a8211d66617c4b59457133ff56fec97f1be591809f187a9f23d04aef670033bc617397df689089271d711b742e6e6de4ab4428287972e600ba0b34edd640f0b5284006ac6c15ea13eb1009e75bc11a0c346e25bbe203e9e7feb1593d7141fdb416e6f26fe8f0d83f2bbe324331c2edbad8f89632d37796fc2a7a8420d4e1d63a3c05e6a4cd58ea468bb7b8950addd10d7eb2588a0e500aed7b25ffa69035fa18e0ec2921387c152782185ec5c90ffe8fc92884d4136ef0ca25119093cbf4ccca232c3943f5873809dd1ddc482eed576f3aa643065313e436feabc6ff139d3ece1b8ccac55a094b23d8a3889171cffbe5872c26515b50d4cff1b1da752052a6a43615617d6d988134a4a8b0c25e74ab44b9941cb88a3b53538aa86b806b1379ea3c7f0bea61f5664dab11abf709dedf91a84577c7099bf03c49e1f6113eda4492272e0467390a89215dc2381b42aef4d276e8378528416f9b53882d56c49a6db8c839ee4d62cb9972f462ed3c7d523a2293170bbb7cd2f26736f785b9e3a23e60154eab20b22f990265bd1f406e082f49ce9f626562fcd1046018d022c3c1428d44185d52be7e73cc72797b6c0e76bbcd61633d526df66a4f242003d31f7a77ba6c5721c55ca8b8b19bc62de148d7aca2486afd0a42401ca4883eb195d0e2308f2bf46446b055f2dccd917f7184b3759cf52d277efa896ca1799304b56d45291803b614be7ec605f9e5381fa18933acc475a86e1c232140d5331ab331557ff370203e8a49478940806eafc461eba12a97903f2c232c4edf1dc7d235b4b7926deee0ac1d8488d09ea3a51245e944ef735fad5122df2808d59db58c7fe0ba4578ef1970f596379e749c5692e2ed61561ba89f0e617fe3df0edba289e728aba67237b8013eeb5c066a332357772f;
    localparam LBP_61 = 10000'ha11beb64f109e664596ec7fb088d3ea30ee217e172aeea4048ebf98188aa9817aec8a8a47eb04577e7a1caa36c8c41c8f2a480e033557b0289ed88b9e1a87af7c3d7a6c33da3006e466071d3a07c09f3541da2319bd04a7d262d957eee4cb8563d4de7974487850e76a487046eb26dab5b6598d166ba66afdc48faaf3a005397778906921ae4b42e71fc50aa82d56af8549136431dd3b3cb442fa97eaf928c305f7d80d5391bb6b4472c11fa76b815febd635130cbeb6660ba517e72eb79e79897ea666cc6212f06ec9868a52c28ed3c8cabdb2a4551b2323ca7a695e1c58940e52cb6ecda0f2d795062ee7610b264741e62d26855b75ed09a764b1a86ce1b675e743df5df02452623ba342700f16009a65883c16fba92c67c820241941a80d6f98f95138bfab2f6b63690dcd405e7aa1cd736283bf58138b94d0a077a0f7a662748c5d2479e01b5890c8468b851ac6887e8fcfdf7f0875ef32118fa536144e79dd1f6c305eddb8b21c1548e007cbedaec8b060e31f7fd96b049bd65126c804dc0ce483a8c93d69430ceb8311bc1f6caef9e6a11b6f50b73794fb285a8d0ecaf21f25b460c36611f400576bd393a5a9b5df09a65e612c8445e66d31257945990cfdb283ef8cab335750b082e06a1377fc074e1a16c84b3a912a5f3968b6568c1c8589fd11bbbd1a7bd219de0d8054cb759fc8b101a5bc1a1fde020931f3a31b0022cc8d9758a300092637a40144ae6b8b01cd6fd6a60bfdcc58e92dfe531fc4d0d66f922671d63399e46bd538e8786b2f2e44fac0d5334d1285a819fa31d1657694487c54510560f81f4a31c459769df2adce0993ce941e7febf128447d5fa5f09002e727470a61e30354cd585d99b9cb44b37aa33adb03f0ff1b6b866e04fabf18231f2e14db669c9b30b5e03ff7f0d464b22d16ac100a65e80195ac91373a0db397b83e605d79779ef7851e783c218fed0e1e1a42ffaa0e451cd42c01ad8f2943a5978e5b685b8216716e96d9da6dc314ed13ac23b3ec300251831bd77f164b750d182fd7097bbcb03205d050a5568df018a55bc3b8d4ec94f1471317301d9630d2eb96a65cd350ef6ef469ecc9964a341f6a6a36ef88068345b21ec038d22af254075a36e9adbf9c4183b8c5fa8107d727e281ca3663e1757ce98273a69dd318edd0215fe38e85f5cdd32a554455e704092ba4f522f1959777ec871e2800bc696a207efaedfeeb2de8f89918b6b5abf32765cf1e8a4a7f8fb78b03d1cae0e57420cade3eaf75e574a1d2c0a3bc94a576a56b523a5a1514df5b1e7b5fc4a32a64c3f08c49d836ddb7b1b19ef11b5a07a045050967dee807437b248244521b9f76a673b2b8a4cbe449cb084f6f7d0c464119ab8c451671847f4cdf50b457286f56dbdb7d2cacc27a44fcd9fb7ae186c0f3bbff119d0e881cdac4cc7475e9ea49bc7d91df00fd71737f7d7b4987a20b1965f24a1ddc8648999d1beb5b1d5cb059e3a0aaf8955bc847b2fe68d9557f4442eddfa773e8add3cfef7ad3384a5ff90e16b61869e69a8c6b03cf61d7cf0ebe8ee9251ab637b3bd5cfec916b68a0884cf1284e157281ad543eb7e32de8d59a3cb6494c9fe3d14cc0cae5ba2ac9aba48c619fee94feede286e9291d58e9711c808038d112e52bf1faaa8c96a5e28ac6933afbdcc2ad5946015fcc642c9d709e114ac2d0b3d5f9109b6ad8b9c1a156bdce176dd6ab06d1ad60f3afe55efb83ee94e485c603c5ea22442cd863f47ffceec128a3;
    localparam LBP_62 = 10000'h14c891535462b2111dc06d99b811a02f13a0741331e029895eda21b5c941232684ed97d27f3611a4b54a3df850af808ce5c0960ddebd5860d30b14eb8527f2cb435422d84c5eec79f4cbd4a1fbf8ce48866e07a97bddb752186e0f8f8b3b1abe8e93a40545f76753b065c98356f68241397c54ba089f4f3bb07cd8c8113dcf23a0ef8f0b31fcc8468cd93b9bacd76bbc18637a4ffc7c9c12bfd1aff198e11e593f68759d80fd08f1bc1eae74a68abb09715efac5fcc938700c55c9a1cf4e8e53fca786e036c3552d024843ff609bf0e993402610aa6ac81466ade6535061d9658cc3742ed3757092d43c0b47809e8c69975cb98db166ad840891d676d5994d8993432018b403ef204c7bfd90561988c59aea50423e1405d33e75c6193f91434d643313a5cbc15c91cd9d33eea84b620c5453847c515fb6c84f1b7a6848d17c2c87d42c38ec9e823c77407d5f74ecca58a2a27073ecd90fbe9c66a0e97862c55a53e8af04a4b6d9cce1141ccd2ea0c0286230a40be1a12b9cc0bf8bd6b4f9ff0c32c96afba8c46ec539a6192990d1cc5e4a7f8a54f52aa93452d68b5a46aec1ca5808ba382f7421a66c886346b47b9aa1a44d04bf3cf059ca979bce4aa68e026d19572c5c4ac0e16749d5d5baa377c9aea1077d2d6cd14259f37e93c9b90953cf2120f61aa82cf5382ae5a62ea7cfdab1aea1dcff0b3baa5fb13545d168410c60be56c79b5095d63cdb0feaba93f6b804184df11c227f6b317fbdbccbc948bc4965b03f3ca65f3b99133060bced1fd162707c26200d8431586bfb0ee9edcbff62d682e843d06463a156880b73c0379158cfc58a1d59687a0be75cef098b1fbb7fcd74fbb30d12f6ad1c97d587c2cd2b46317d289f714a0a001554bb1ea2deb3132c06c7b9e405650049fcd5db431fc7d4c5a51251ba3c2cf346259fddfbbccf1db7cc96a3ede920051e87b350a0ddd54b7f95e6196a0c473b6099a18da45ca84d27e69630ed29ff40e3b98a125514ed435e01965c0f0a7652fad0f1c985ed0ae2035adaed0773e4dc6995079a32c7d50e2b5a7db95755e5c3b16542b7f7b2fc0076da9f83ef7da5fe9dbdf776e3e688ec4c13d69fa15eb01745e809af163353e43d7af5897534d7065443d30c67815a0cee627659259c60a5c66adae5456d7da712c60875f021b88c99f5f7c5a052d69cb3cf74d6cdc0174fcff9d3ca666647d2e0c3a33a6c602d743c14a28d40fbcc05895a7f3991968dc2b30ebff6420cb99c3228dfc7d5e9b4c4ec130e4a934afbc16c7c793bb3af5e1716cccb7d3298e8c8811a72fc359c44937e411159f0fa8169ab3024965497b642ead4ffb4d600c0a6e72c0a4a7a4e8ecd69f5ab2f1951a817470e0e140edeb236341d337605a12f27a0526af88a6e21fb0dfe947c23ec76847b40bb003aa86fdb9bf53bf5ef71a94a85fb04762dcda43a94cad974798f4663fb94b67ebf9d428a5702ea29e27d75a1ceed71f17cf705955ce44e2fcfc8ebe706f0956fd6d565f6ff38bc08efe503e4b5689058d9cddeddbd3f7acb9699a5235a90aec41ba44b285b7319866350dff39b52d212123bb5c598d998cb926ee12db00e89c08034ad7cfa9cc62adce17430e543d93f2f8068df025c52b012463108b5032e10b211e070e71307f23c25b5a465ae725583e6852b21bf6ef7d444cd08c2df57808725f3f4feb2a8783b34fed277cce283de9b85274b63feb428065d99908f0244fc83a26da13daa628af7b272afdd;
    localparam LBP_63 = 10000'hd5801c873bbed0a0d7aa3bc74eaa2731689549ae1ce7052969a13c07f28f2664e445551a8635591f316960521db424403abf957cf71cd54adeb35c5147e0e7c62f5544234b0338e9684180cd329ab9c93893ed25cb3fbfd55833f30feaf2bdb669c4c5cff7550eb64aaf59598272a933a538b927941fec799c717909d880a42379537349fe78e4141200e1d5f1f065529e0bdf73864d105c5a34c21448d737d8282a90ab10ad383872cdd64a0497a22aa5bf51e89ff4b1d73b7a0acb14c2617ac95a7c346176bbff4cf0a2ec93f007748b3f80781727c2d5531e1130b49a9d1709e97d6e5ad172d3c82debdf7748606def7bf6a258532bd664c1f4ec7478629a50e95151c90a705a816205bdb15dd1263d96f2c7b44153448817420534f7de13e36a6e681912add308bd8c19ca0f8e4ad7d3ea218508b9df7b898186cc1d1a8cbd2070d31fdd4bbddc62d42ca93231e4f0079600904219c1ba261e47e59db70b90f02693ed622d3204b3182001c0410823692f2ef50d38123d1f5025076ef0aa592ccb2dc930b9727345d63f3d62abe80bca9f93c16c34686166652159aa0b73c23fd3dc441712ae328eae92e7def6ad6aefe4e760b5daa0f32fa0ceaf249809836f6a04fd1b44076f649fde92a7b473f57d3008090871cc9fe6fdb6bfb7c09d76efd224bbecfff2e41442f8528866d48616f924f9c910a026ddc7f33a3d316d3e8d8ba6a164307af3207b842a3fdc52f69b438c828c9668d7d11b4ac8bed345c3fc8b02dcba619d5341d19a884792ffc0e07fe2702820144fd1f948edf683e83190fd245d65d8e4854dbbebab0834aae7420056fff434a429837f59dff429a1d20ce0c2f1954753eb7d5502855c58a66bd879996afa6a480a14cdf5d4340edb36ccf5d1691e7565679b81e90bf346caadfade3183a6bfac3f57d7f1ddc73b113ef0d11a5636a1fa68ec0c258c58946cb573db5a8ccce19698669aa50886fe0335fe7845b9c400859000f9385a4d1c3c46a46a9aa5f22b039eb34a52325afa996f921d41ad3c1f3d860afc69ca6cf93746c118a841f39da7c7803af5a0f15c2fecd2c995c39b70ec5f68e10c65775b3cca6375b3e2c9f1a0ecf4d2db84fceacb11fd798bc1d2c46dec43fd6d81ccb76bbba2da3f8a7b5b68efb9a1fbdb1092e36bc37b39d401a85ed6bc623fa3f57015f358874fead3a2070e77f8bcbeb73a08f9c2d2e9c67639f8daf55a2c5910c5338077865f2d5be28b83f9d5f8efadf105266ef4fa6bdd4043c25544102f2d6b3026593053a39209153b0de63ff1643c8daaf7e1a11532ff7fa84c997789217d7fdac45fce2b917397f095aeefe312a39ccc32c0259b86135c85c138a603d3f1e5ed197f418f4754e03510d1dce90a6376f707cc53ea4ed41c4d063eea820018c5ea95864353663587b6f9adaa0ae59a3586597264838970b262808ffb8ffedbaca0ca76b070216f5a855e007758a8a0cff3f2d43b59c97938db6921d07c3441817dc59892a67420250d62388098726a8c8b53427f4daba38c24d295603f9f4559a694fae0b187cec112b7323fc0bf2fb8e49a31908c7fdd3a4dfde733d19d4ada3e78897a3a5348677ae56783ecb757320b9626f419835d388e2b2948ecee40e0209707f59362ebedeaddc25eee258269561b9430c8cdf54b2d3438eb6cd1bb7f250ec9a56897cb5c8d0b8443c55f1c6b438f6b7b4bd014da73dea682aaf5d349114a2262f68f8c8af37eaea4b719593236fd;


    input [$clog2(NUM_CHS) - 1: 0] c;
    input [$clog2(NUM_LBP) - 1: 0] l;
    output logic [DIMENSIONS - 1:0] ch_hv;
    output logic [DIMENSIONS - 1:0] lbp_hv;


    wire [NUM_CHS - 1: 0][DIMENSIONS - 1:0] ch_mem;
    wire [NUM_LBP - 1: 0][DIMENSIONS - 1:0] lbp_mem;


    assign ch_mem[0] = CH_0;
    assign ch_mem[1] = CH_1;
    assign ch_mem[2] = CH_2;
    assign ch_mem[3] = CH_3;
    assign ch_mem[4] = CH_4;
    assign ch_mem[5] = CH_5;
    assign ch_mem[6] = CH_6;
    assign ch_mem[7] = CH_7;
    assign ch_mem[8] = CH_8;
    assign ch_mem[9] = CH_9;
    assign ch_mem[10] = CH_10;
    assign ch_mem[11] = CH_11;
    assign ch_mem[12] = CH_12;
    assign ch_mem[13] = CH_13;
    assign ch_mem[14] = CH_14;
    assign ch_mem[15] = CH_15;
    assign ch_mem[16] = CH_16;


    assign lbp_mem[0] = LBP_0;
    assign lbp_mem[1] = LBP_1;
    assign lbp_mem[2] = LBP_2;
    assign lbp_mem[3] = LBP_3;
    assign lbp_mem[4] = LBP_4;
    assign lbp_mem[5] = LBP_5;
    assign lbp_mem[6] = LBP_6;
    assign lbp_mem[7] = LBP_7;
    assign lbp_mem[8] = LBP_8;
    assign lbp_mem[9] = LBP_9;
    assign lbp_mem[10] = LBP_10;
    assign lbp_mem[11] = LBP_11;
    assign lbp_mem[12] = LBP_12;
    assign lbp_mem[13] = LBP_13;
    assign lbp_mem[14] = LBP_14;
    assign lbp_mem[15] = LBP_15;
    assign lbp_mem[16] = LBP_16;
    assign lbp_mem[17] = LBP_17;
    assign lbp_mem[18] = LBP_18;
    assign lbp_mem[19] = LBP_19;
    assign lbp_mem[20] = LBP_20;
    assign lbp_mem[21] = LBP_21;
    assign lbp_mem[22] = LBP_22;
    assign lbp_mem[23] = LBP_23;
    assign lbp_mem[24] = LBP_24;
    assign lbp_mem[25] = LBP_25;
    assign lbp_mem[26] = LBP_26;
    assign lbp_mem[27] = LBP_27;
    assign lbp_mem[28] = LBP_28;
    assign lbp_mem[29] = LBP_29;
    assign lbp_mem[30] = LBP_30;
    assign lbp_mem[31] = LBP_31;
    assign lbp_mem[32] = LBP_32;
    assign lbp_mem[33] = LBP_33;
    assign lbp_mem[34] = LBP_34;
    assign lbp_mem[35] = LBP_35;
    assign lbp_mem[36] = LBP_36;
    assign lbp_mem[37] = LBP_37;
    assign lbp_mem[38] = LBP_38;
    assign lbp_mem[39] = LBP_39;
    assign lbp_mem[40] = LBP_40;
    assign lbp_mem[41] = LBP_41;
    assign lbp_mem[42] = LBP_42;
    assign lbp_mem[43] = LBP_43;
    assign lbp_mem[44] = LBP_44;
    assign lbp_mem[45] = LBP_45;
    assign lbp_mem[46] = LBP_46;
    assign lbp_mem[47] = LBP_47;
    assign lbp_mem[48] = LBP_48;
    assign lbp_mem[49] = LBP_49;
    assign lbp_mem[50] = LBP_50;
    assign lbp_mem[51] = LBP_51;
    assign lbp_mem[52] = LBP_52;
    assign lbp_mem[53] = LBP_53;
    assign lbp_mem[54] = LBP_54;
    assign lbp_mem[55] = LBP_55;
    assign lbp_mem[56] = LBP_56;
    assign lbp_mem[57] = LBP_57;
    assign lbp_mem[58] = LBP_58;
    assign lbp_mem[59] = LBP_59;
    assign lbp_mem[60] = LBP_60;
    assign lbp_mem[61] = LBP_61;
    assign lbp_mem[62] = LBP_62;
    assign lbp_mem[63] = LBP_63;

    always_comb begin
        ch_hv = ch_mem[c];
        lbp_hv = lbp_mem[l];
    end

endmodule