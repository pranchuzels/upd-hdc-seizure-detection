`timescale 1us / 1ns
module tb_ma_encoder_mapped ();
    localparam T = 1.0;  // clock period in us

    // General params
    localparam DIMENSIONS = 10000;
    localparam NUM_CHS = 17;
    localparam WINDOW_SIZE = 256;
    localparam WINDOW_STEP = 128;
    localparam SAMPLE_SIZE = 16;

    // Feature params
    parameter NUM_MA = 64;

    // Bundler params
    localparam COUNT_SIZE = 8;

    reg clk;
    reg nrst;
    reg en;
    reg [NUM_CHS - 1: 0][SAMPLE_SIZE - 1: 0] samples;
    wire done;
    wire [DIMENSIONS - 1:0] window_hv;

    ma_encoder #(
        .DIMENSIONS(DIMENSIONS),
        .NUM_CHS(NUM_CHS),
        .WINDOW_SIZE(WINDOW_SIZE),
        .WINDOW_STEP(WINDOW_STEP),
        .SAMPLE_SIZE(SAMPLE_SIZE),
        .NUM_MA(NUM_MA),
        .COUNT_SIZE(COUNT_SIZE)
    )
    u_ma_encoder(   
        .clk (clk),
        .nrst (nrst),
        .en (en),
        .samples (samples),
        .done (done),
        .window_hv (window_hv)
    );

    // Clock
    always begin
        clk = 1'b1;
        #(T / 2.0);
        clk = 1'b0;
        #(T / 2.0);

        if ($time % 100000 == 0) begin
            $display("Current time is: %t", $time);
        end
        //$display("Current time is: %t", $time);
    end

    initial begin
        $sdf_annotate("../mapped/ma_encoder_mapped.sdf", u_ma_encoder);

        nrst = 0;
        en = 0;
        samples = 0;
        # (10 - 0.5)
        nrst = 1;

        en = 1;
        samples[0] = 16'b1111110111101011;
        samples[1] = 16'b1111111101010110;
        samples[2] = 16'b1111110111110100;
        samples[3] = 16'b1111111110100001;
        samples[4] = 16'b1111110111001001;
        samples[5] = 16'b1111111001110001;
        samples[6] = 16'b1111111010110011;
        samples[7] = 16'b1111111111101100;
        samples[8] = 16'b1111110111111110;
        samples[9] = 16'b1111110100101100;
        samples[10] = 16'b1111111101001100;
        samples[11] = 16'b1111111010010111;
        samples[12] = 16'b1111101001100111;
        samples[13] = 16'b1111110110001010;
        samples[14] = 16'b1111111010101101;
        samples[15] = 16'b1111110110000100;
        samples[16] = 16'b1111111101010110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111000111001;
        samples[1] = 16'b1111111101111000;
        samples[2] = 16'b1111111000000111;
        samples[3] = 16'b1111111101011001;
        samples[4] = 16'b1111111000000001;
        samples[5] = 16'b1111111010010111;
        samples[6] = 16'b1111111011001111;
        samples[7] = 16'b1111111110100111;
        samples[8] = 16'b1111111010001110;
        samples[9] = 16'b1111110010010110;
        samples[10] = 16'b1111111101001100;
        samples[11] = 16'b1111111100000100;
        samples[12] = 16'b1111110000111100;
        samples[13] = 16'b1111110100101001;
        samples[14] = 16'b1111111100100111;
        samples[15] = 16'b1111110110001010;
        samples[16] = 16'b1111111100111010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111001110101;
        samples[1] = 16'b1111111110000001;
        samples[2] = 16'b1111111000000001;
        samples[3] = 16'b1111111101101111;
        samples[4] = 16'b1111111001000011;
        samples[5] = 16'b1111111010011010;
        samples[6] = 16'b1111111011001100;
        samples[7] = 16'b1111111110111010;
        samples[8] = 16'b1111111000111100;
        samples[9] = 16'b1111110100101001;
        samples[10] = 16'b1111111100111010;
        samples[11] = 16'b1111111101000110;
        samples[12] = 16'b1111110110110011;
        samples[13] = 16'b1111110001111010;
        samples[14] = 16'b1111111110000101;
        samples[15] = 16'b1111110111001001;
        samples[16] = 16'b1111111100001011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011001111;
        samples[1] = 16'b1111111110110011;
        samples[2] = 16'b1111111000101010;
        samples[3] = 16'b1111111100111101;
        samples[4] = 16'b1111111010100111;
        samples[5] = 16'b1111111010110000;
        samples[6] = 16'b1111111011001001;
        samples[7] = 16'b1111111111001001;
        samples[8] = 16'b1111111001001100;
        samples[9] = 16'b1111110110011010;
        samples[10] = 16'b1111111101001100;
        samples[11] = 16'b1111111100011010;
        samples[12] = 16'b1111110100001101;
        samples[13] = 16'b1111111101011100;
        samples[14] = 16'b1111111010101101;
        samples[15] = 16'b1111110111111110;
        samples[16] = 16'b1111111011101011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100100100;
        samples[1] = 16'b1111111111011001;
        samples[2] = 16'b1111111000111100;
        samples[3] = 16'b1111111100000001;
        samples[4] = 16'b1111111011111011;
        samples[5] = 16'b1111111010101010;
        samples[6] = 16'b1111111010111100;
        samples[7] = 16'b1111111111010110;
        samples[8] = 16'b1111111010111001;
        samples[9] = 16'b1111110100111100;
        samples[10] = 16'b1111111101001001;
        samples[11] = 16'b1111111110001011;
        samples[12] = 16'b1111110011111101;
        samples[13] = 16'b1111110111111110;
        samples[14] = 16'b1111111100100111;
        samples[15] = 16'b1111111000001101;
        samples[16] = 16'b1111111010110011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101110010;
        samples[1] = 16'b1111111111000000;
        samples[2] = 16'b1111111001010010;
        samples[3] = 16'b1111111011110010;
        samples[4] = 16'b1111111100100111;
        samples[5] = 16'b1111111010001110;
        samples[6] = 16'b1111111011000011;
        samples[7] = 16'b1111111111111011;
        samples[8] = 16'b1111111000000001;
        samples[9] = 16'b1111110110001101;
        samples[10] = 16'b1111111111010000;
        samples[11] = 16'b1111111111101001;
        samples[12] = 16'b1111110100011101;
        samples[13] = 16'b1111110100110000;
        samples[14] = 16'b1111111101001001;
        samples[15] = 16'b1111111000111100;
        samples[16] = 16'b1111111010100111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110100111;
        samples[1] = 16'b1111111110100100;
        samples[2] = 16'b1111111001101011;
        samples[3] = 16'b1111111010110011;
        samples[4] = 16'b1111111100111010;
        samples[5] = 16'b1111111001101110;
        samples[6] = 16'b1111111010100000;
        samples[7] = 16'b0000000000011011;
        samples[8] = 16'b1111110110000001;
        samples[9] = 16'b1111110110110000;
        samples[10] = 16'b0000000000100111;
        samples[11] = 16'b1111111101101100;
        samples[12] = 16'b1111110011101011;
        samples[13] = 16'b1111111101000110;
        samples[14] = 16'b1111111011000110;
        samples[15] = 16'b1111111000111100;
        samples[16] = 16'b1111111001111000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110100111;
        samples[1] = 16'b1111111101111011;
        samples[2] = 16'b1111111001011100;
        samples[3] = 16'b1111111010101101;
        samples[4] = 16'b1111111100100111;
        samples[5] = 16'b1111111000110011;
        samples[6] = 16'b1111111001110101;
        samples[7] = 16'b0000000001011100;
        samples[8] = 16'b1111110100101001;
        samples[9] = 16'b1111110111111011;
        samples[10] = 16'b0000000000001000;
        samples[11] = 16'b1111111100011101;
        samples[12] = 16'b1111110001001110;
        samples[13] = 16'b0000000011101111;
        samples[14] = 16'b1111111010010111;
        samples[15] = 16'b1111111000111001;
        samples[16] = 16'b1111111001000011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111111010011;
        samples[1] = 16'b1111111100111010;
        samples[2] = 16'b1111111001111110;
        samples[3] = 16'b1111111010110000;
        samples[4] = 16'b1111111101010011;
        samples[5] = 16'b1111111000001010;
        samples[6] = 16'b1111111010010100;
        samples[7] = 16'b0000000001000011;
        samples[8] = 16'b1111110101100010;
        samples[9] = 16'b1111111010011010;
        samples[10] = 16'b1111111110001110;
        samples[11] = 16'b1111111101010011;
        samples[12] = 16'b1111110011001011;
        samples[13] = 16'b0000000001100110;
        samples[14] = 16'b1111111100001011;
        samples[15] = 16'b1111111001101011;
        samples[16] = 16'b1111111001100101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111111000110;
        samples[1] = 16'b1111111011110010;
        samples[2] = 16'b1111111001111000;
        samples[3] = 16'b1111111100001011;
        samples[4] = 16'b1111111101001111;
        samples[5] = 16'b1111110110101101;
        samples[6] = 16'b1111111010101010;
        samples[7] = 16'b0000000010010001;
        samples[8] = 16'b1111110100010000;
        samples[9] = 16'b1111111011000110;
        samples[10] = 16'b1111111110000001;
        samples[11] = 16'b1111111110001110;
        samples[12] = 16'b1111111010011010;
        samples[13] = 16'b0000001010011000;
        samples[14] = 16'b1111111101000110;
        samples[15] = 16'b1111111001111110;
        samples[16] = 16'b1111111001111000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101000011;
        samples[1] = 16'b1111111010111100;
        samples[2] = 16'b1111111010000100;
        samples[3] = 16'b1111111110110111;
        samples[4] = 16'b1111111011011111;
        samples[5] = 16'b1111110100110000;
        samples[6] = 16'b1111111010010111;
        samples[7] = 16'b0000000110010010;
        samples[8] = 16'b1111110011001111;
        samples[9] = 16'b1111111101000110;
        samples[10] = 16'b1111111011101110;
        samples[11] = 16'b1111111101110101;
        samples[12] = 16'b1111110110111111;
        samples[13] = 16'b0000000101110110;
        samples[14] = 16'b1111111001101000;
        samples[15] = 16'b1111111010000100;
        samples[16] = 16'b1111111000111100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101000110;
        samples[1] = 16'b1111111011010101;
        samples[2] = 16'b1111111010100000;
        samples[3] = 16'b1111111110001011;
        samples[4] = 16'b1111111011011100;
        samples[5] = 16'b1111110100111100;
        samples[6] = 16'b1111111011001100;
        samples[7] = 16'b0000000101100000;
        samples[8] = 16'b1111110011010010;
        samples[9] = 16'b1111111100100100;
        samples[10] = 16'b1111111100110011;
        samples[11] = 16'b1111111101100010;
        samples[12] = 16'b1111111001000110;
        samples[13] = 16'b0000000110011110;
        samples[14] = 16'b1111111001011100;
        samples[15] = 16'b1111111010111001;
        samples[16] = 16'b1111111001111110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101000011;
        samples[1] = 16'b1111111010110000;
        samples[2] = 16'b1111111011001100;
        samples[3] = 16'b1111111110101010;
        samples[4] = 16'b1111111011000011;
        samples[5] = 16'b1111110100110110;
        samples[6] = 16'b1111111100100111;
        samples[7] = 16'b0000000101000100;
        samples[8] = 16'b1111110000100110;
        samples[9] = 16'b1111111011100010;
        samples[10] = 16'b1111111111111110;
        samples[11] = 16'b1111111110010100;
        samples[12] = 16'b1111111100100001;
        samples[13] = 16'b0000000010101101;
        samples[14] = 16'b1111111011111110;
        samples[15] = 16'b1111111011010101;
        samples[16] = 16'b1111111011001111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101100010;
        samples[1] = 16'b1111111010110011;
        samples[2] = 16'b1111111011101000;
        samples[3] = 16'b1111111101110101;
        samples[4] = 16'b1111111011100010;
        samples[5] = 16'b1111110110100110;
        samples[6] = 16'b1111111100110110;
        samples[7] = 16'b0000000010110001;
        samples[8] = 16'b1111110011011110;
        samples[9] = 16'b1111111100100100;
        samples[10] = 16'b1111111111010011;
        samples[11] = 16'b1111111011101110;
        samples[12] = 16'b1111111011101011;
        samples[13] = 16'b0000000110011110;
        samples[14] = 16'b1111111011101110;
        samples[15] = 16'b1111111011110101;
        samples[16] = 16'b1111111011001100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101101000;
        samples[1] = 16'b1111111010101010;
        samples[2] = 16'b1111111100001000;
        samples[3] = 16'b1111111101011111;
        samples[4] = 16'b1111111011110010;
        samples[5] = 16'b1111111000000001;
        samples[6] = 16'b1111111100101010;
        samples[7] = 16'b0000000001010110;
        samples[8] = 16'b1111110110010000;
        samples[9] = 16'b1111111101000110;
        samples[10] = 16'b1111111101111000;
        samples[11] = 16'b1111111010111001;
        samples[12] = 16'b1111111100100001;
        samples[13] = 16'b1111111111000011;
        samples[14] = 16'b1111111001111110;
        samples[15] = 16'b1111111100000001;
        samples[16] = 16'b1111111011010010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101111110;
        samples[1] = 16'b1111111010100011;
        samples[2] = 16'b1111111100011010;
        samples[3] = 16'b1111111101011001;
        samples[4] = 16'b1111111100011101;
        samples[5] = 16'b1111111001001100;
        samples[6] = 16'b1111111100110011;
        samples[7] = 16'b1111111111101111;
        samples[8] = 16'b1111111011111000;
        samples[9] = 16'b1111111111110101;
        samples[10] = 16'b1111111001101110;
        samples[11] = 16'b1111111000100000;
        samples[12] = 16'b1111111110011110;
        samples[13] = 16'b0000000010101010;
        samples[14] = 16'b1111110111101011;
        samples[15] = 16'b1111111100101010;
        samples[16] = 16'b1111111011010010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101010011;
        samples[1] = 16'b1111111010000100;
        samples[2] = 16'b1111111100001000;
        samples[3] = 16'b1111111110110000;
        samples[4] = 16'b1111111011110101;
        samples[5] = 16'b1111111001001111;
        samples[6] = 16'b1111111101000000;
        samples[7] = 16'b0000000000000010;
        samples[8] = 16'b1111111011101011;
        samples[9] = 16'b1111111111111000;
        samples[10] = 16'b1111111010011101;
        samples[11] = 16'b1111110111110001;
        samples[12] = 16'b0000000100001000;
        samples[13] = 16'b1111111110010100;
        samples[14] = 16'b1111110101001001;
        samples[15] = 16'b1111111100111101;
        samples[16] = 16'b1111111010110110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101000011;
        samples[1] = 16'b1111111010011101;
        samples[2] = 16'b1111111101001001;
        samples[3] = 16'b1111111110100111;
        samples[4] = 16'b1111111011101011;
        samples[5] = 16'b1111111001110001;
        samples[6] = 16'b1111111101111011;
        samples[7] = 16'b1111111111110010;
        samples[8] = 16'b1111111101000000;
        samples[9] = 16'b0000000010010001;
        samples[10] = 16'b1111111001011111;
        samples[11] = 16'b1111110111000110;
        samples[12] = 16'b0000000011011100;
        samples[13] = 16'b1111111110011110;
        samples[14] = 16'b1111110011110100;
        samples[15] = 16'b1111111101100101;
        samples[16] = 16'b1111111011000000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101001111;
        samples[1] = 16'b1111111010101101;
        samples[2] = 16'b1111111101011111;
        samples[3] = 16'b1111111110100001;
        samples[4] = 16'b1111111011110101;
        samples[5] = 16'b1111111010000100;
        samples[6] = 16'b1111111110011010;
        samples[7] = 16'b1111111111101100;
        samples[8] = 16'b1111111110100001;
        samples[9] = 16'b0000000000000010;
        samples[10] = 16'b1111111001111011;
        samples[11] = 16'b1111111000010100;
        samples[12] = 16'b0000000010110111;
        samples[13] = 16'b1111111110000101;
        samples[14] = 16'b1111110110000001;
        samples[15] = 16'b1111111101100010;
        samples[16] = 16'b1111111011011100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101011001;
        samples[1] = 16'b1111111011011001;
        samples[2] = 16'b1111111101111110;
        samples[3] = 16'b1111111101001100;
        samples[4] = 16'b1111111011110101;
        samples[5] = 16'b1111111010100011;
        samples[6] = 16'b1111111111000110;
        samples[7] = 16'b1111111110011110;
        samples[8] = 16'b1111111101011100;
        samples[9] = 16'b1111111101000011;
        samples[10] = 16'b1111111100010111;
        samples[11] = 16'b1111111000010100;
        samples[12] = 16'b1111111111011100;
        samples[13] = 16'b1111111100101010;
        samples[14] = 16'b1111110111010101;
        samples[15] = 16'b1111111100101101;
        samples[16] = 16'b1111111100000100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101011111;
        samples[1] = 16'b1111111100001000;
        samples[2] = 16'b1111111110100111;
        samples[3] = 16'b1111111100101010;
        samples[4] = 16'b1111111100011010;
        samples[5] = 16'b1111111011001111;
        samples[6] = 16'b1111111111011100;
        samples[7] = 16'b1111111101110101;
        samples[8] = 16'b1111111111001100;
        samples[9] = 16'b1111111101101100;
        samples[10] = 16'b1111111010100111;
        samples[11] = 16'b1111111000001101;
        samples[12] = 16'b1111110110101101;
        samples[13] = 16'b0000000110110111;
        samples[14] = 16'b1111111000010001;
        samples[15] = 16'b1111111100011101;
        samples[16] = 16'b1111111100011101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101101000;
        samples[1] = 16'b1111111100001000;
        samples[2] = 16'b1111111110011010;
        samples[3] = 16'b1111111100101010;
        samples[4] = 16'b1111111101001001;
        samples[5] = 16'b1111111011010010;
        samples[6] = 16'b1111111111011001;
        samples[7] = 16'b1111111100111010;
        samples[8] = 16'b0000000000001000;
        samples[9] = 16'b1111111101011001;
        samples[10] = 16'b1111111001011111;
        samples[11] = 16'b1111111010010111;
        samples[12] = 16'b1111111010110011;
        samples[13] = 16'b1111111100011101;
        samples[14] = 16'b1111111010011010;
        samples[15] = 16'b1111111100001110;
        samples[16] = 16'b1111111101000110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110010111;
        samples[1] = 16'b1111111100101101;
        samples[2] = 16'b1111111110011010;
        samples[3] = 16'b1111111011101110;
        samples[4] = 16'b1111111110100001;
        samples[5] = 16'b1111111011011001;
        samples[6] = 16'b0000000000000010;
        samples[7] = 16'b1111111011000110;
        samples[8] = 16'b1111111111011111;
        samples[9] = 16'b1111111101011100;
        samples[10] = 16'b1111111011011111;
        samples[11] = 16'b1111111100011010;
        samples[12] = 16'b1111111101000000;
        samples[13] = 16'b1111111111101100;
        samples[14] = 16'b1111111100001011;
        samples[15] = 16'b1111111100001110;
        samples[16] = 16'b1111111110001110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110001000;
        samples[1] = 16'b1111111101000110;
        samples[2] = 16'b1111111110001011;
        samples[3] = 16'b1111111011110101;
        samples[4] = 16'b1111111110110000;
        samples[5] = 16'b1111111010100000;
        samples[6] = 16'b1111111111111011;
        samples[7] = 16'b1111111011110010;
        samples[8] = 16'b1111111100010100;
        samples[9] = 16'b1111111100100001;
        samples[10] = 16'b1111111101011001;
        samples[11] = 16'b1111111110001011;
        samples[12] = 16'b1111111100000001;
        samples[13] = 16'b0000000110111010;
        samples[14] = 16'b1111111110010111;
        samples[15] = 16'b1111111011100101;
        samples[16] = 16'b1111111110010001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101010011;
        samples[1] = 16'b1111111101000000;
        samples[2] = 16'b1111111101101111;
        samples[3] = 16'b1111111100010100;
        samples[4] = 16'b1111111110011110;
        samples[5] = 16'b1111111000111100;
        samples[6] = 16'b1111111111110010;
        samples[7] = 16'b1111111101000011;
        samples[8] = 16'b1111111001100101;
        samples[9] = 16'b1111111011000011;
        samples[10] = 16'b1111111110110000;
        samples[11] = 16'b0000000000100100;
        samples[12] = 16'b1111111111100101;
        samples[13] = 16'b1111110000101001;
        samples[14] = 16'b1111111111111000;
        samples[15] = 16'b1111111010111001;
        samples[16] = 16'b1111111110100100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101001001;
        samples[1] = 16'b1111111011111000;
        samples[2] = 16'b1111111101001100;
        samples[3] = 16'b1111111100110110;
        samples[4] = 16'b1111111101111000;
        samples[5] = 16'b1111110111001111;
        samples[6] = 16'b0000000000101010;
        samples[7] = 16'b1111111101001001;
        samples[8] = 16'b1111110111111011;
        samples[9] = 16'b1111111010000100;
        samples[10] = 16'b0000000000011011;
        samples[11] = 16'b0000000100000101;
        samples[12] = 16'b1111111101100010;
        samples[13] = 16'b1111110100100110;
        samples[14] = 16'b0000000101011001;
        samples[15] = 16'b1111111010010111;
        samples[16] = 16'b1111111111110010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011101110;
        samples[1] = 16'b1111111010100011;
        samples[2] = 16'b1111111101001001;
        samples[3] = 16'b1111111110000001;
        samples[4] = 16'b1111111100011101;
        samples[5] = 16'b1111110101000010;
        samples[6] = 16'b0000000001010000;
        samples[7] = 16'b1111111110011110;
        samples[8] = 16'b1111111000001010;
        samples[9] = 16'b1111111000111100;
        samples[10] = 16'b1111111110101101;
        samples[11] = 16'b0000000111001010;
        samples[12] = 16'b1111110110111100;
        samples[13] = 16'b1111111000000111;
        samples[14] = 16'b0000001001010111;
        samples[15] = 16'b1111111001000011;
        samples[16] = 16'b0000000000000010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111010100000;
        samples[1] = 16'b1111111010100000;
        samples[2] = 16'b1111111100111010;
        samples[3] = 16'b1111111110101101;
        samples[4] = 16'b1111111010101010;
        samples[5] = 16'b1111110100101001;
        samples[6] = 16'b0000000001001001;
        samples[7] = 16'b0000000000000010;
        samples[8] = 16'b1111110101110111;
        samples[9] = 16'b1111111010101010;
        samples[10] = 16'b1111111111100101;
        samples[11] = 16'b0000000110110100;
        samples[12] = 16'b1111110001101110;
        samples[13] = 16'b1111101010111110;
        samples[14] = 16'b0000000110011000;
        samples[15] = 16'b1111111000110110;
        samples[16] = 16'b0000000000110000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111010111001;
        samples[1] = 16'b1111111011110010;
        samples[2] = 16'b1111111101011100;
        samples[3] = 16'b1111111100110000;
        samples[4] = 16'b1111111010010001;
        samples[5] = 16'b1111110110000111;
        samples[6] = 16'b0000000001111011;
        samples[7] = 16'b1111111110010100;
        samples[8] = 16'b1111110111101110;
        samples[9] = 16'b1111111011001111;
        samples[10] = 16'b0000000000100001;
        samples[11] = 16'b0000000101000000;
        samples[12] = 16'b1111110011110111;
        samples[13] = 16'b1111111010011010;
        samples[14] = 16'b0000000101110010;
        samples[15] = 16'b1111111001000110;
        samples[16] = 16'b0000000011001101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011011001;
        samples[1] = 16'b1111111011111011;
        samples[2] = 16'b1111111101000011;
        samples[3] = 16'b1111111101001001;
        samples[4] = 16'b1111111001100101;
        samples[5] = 16'b1111110111110001;
        samples[6] = 16'b0000000010011110;
        samples[7] = 16'b1111111101011100;
        samples[8] = 16'b1111110101111011;
        samples[9] = 16'b1111111101010110;
        samples[10] = 16'b0000000010111101;
        samples[11] = 16'b0000000101111111;
        samples[12] = 16'b1111110000110010;
        samples[13] = 16'b1111110111100101;
        samples[14] = 16'b0000000101101001;
        samples[15] = 16'b1111111001010101;
        samples[16] = 16'b0000000101100000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100100001;
        samples[1] = 16'b1111111101001001;
        samples[2] = 16'b1111111100101101;
        samples[3] = 16'b1111111100001110;
        samples[4] = 16'b1111111001001111;
        samples[5] = 16'b1111111001101011;
        samples[6] = 16'b0000000011000011;
        samples[7] = 16'b1111111100010111;
        samples[8] = 16'b1111110010111111;
        samples[9] = 16'b1111111110100001;
        samples[10] = 16'b0000000110111010;
        samples[11] = 16'b0000000110101000;
        samples[12] = 16'b1111110111010101;
        samples[13] = 16'b1111110110000100;
        samples[14] = 16'b0000000101111100;
        samples[15] = 16'b1111111010011010;
        samples[16] = 16'b0000000111100110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100101010;
        samples[1] = 16'b1111111101010110;
        samples[2] = 16'b1111111011111000;
        samples[3] = 16'b1111111100001011;
        samples[4] = 16'b1111111000000100;
        samples[5] = 16'b1111111010100111;
        samples[6] = 16'b0000000010110111;
        samples[7] = 16'b1111111100010100;
        samples[8] = 16'b1111110011000010;
        samples[9] = 16'b1111111101101111;
        samples[10] = 16'b0000000111010011;
        samples[11] = 16'b0000001000100101;
        samples[12] = 16'b1111111001010010;
        samples[13] = 16'b1111110110011010;
        samples[14] = 16'b0000000111111001;
        samples[15] = 16'b1111111011000011;
        samples[16] = 16'b0000001000100001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100100111;
        samples[1] = 16'b1111111101010110;
        samples[2] = 16'b1111111011010010;
        samples[3] = 16'b1111111101000110;
        samples[4] = 16'b1111110110100011;
        samples[5] = 16'b1111111011001111;
        samples[6] = 16'b0000000011010110;
        samples[7] = 16'b1111111100111101;
        samples[8] = 16'b1111110001001011;
        samples[9] = 16'b1111111110011010;
        samples[10] = 16'b0000001000101000;
        samples[11] = 16'b0000001010011000;
        samples[12] = 16'b1111111001101110;
        samples[13] = 16'b1111111110100001;
        samples[14] = 16'b0000001000101110;
        samples[15] = 16'b1111111100001000;
        samples[16] = 16'b0000001001000111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011010101;
        samples[1] = 16'b1111111101001100;
        samples[2] = 16'b1111111010110110;
        samples[3] = 16'b1111111110100001;
        samples[4] = 16'b1111110100100000;
        samples[5] = 16'b1111111011011001;
        samples[6] = 16'b0000000011101100;
        samples[7] = 16'b1111111101111110;
        samples[8] = 16'b1111110000010000;
        samples[9] = 16'b0000000000100100;
        samples[10] = 16'b0000000111011010;
        samples[11] = 16'b0000001001110011;
        samples[12] = 16'b1111111011011111;
        samples[13] = 16'b1111110101011011;
        samples[14] = 16'b0000001000000101;
        samples[15] = 16'b1111111100110000;
        samples[16] = 16'b0000001001000100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011110101;
        samples[1] = 16'b1111111101111110;
        samples[2] = 16'b1111111010101010;
        samples[3] = 16'b1111111110100100;
        samples[4] = 16'b1111110100000001;
        samples[5] = 16'b1111111100101101;
        samples[6] = 16'b0000000100000010;
        samples[7] = 16'b1111111110000001;
        samples[8] = 16'b1111110010001010;
        samples[9] = 16'b1111111111111110;
        samples[10] = 16'b0000000111111100;
        samples[11] = 16'b0000001010011011;
        samples[12] = 16'b1111110101000010;
        samples[13] = 16'b0000000111000100;
        samples[14] = 16'b0000001000101110;
        samples[15] = 16'b1111111101111000;
        samples[16] = 16'b0000001001010000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100000100;
        samples[1] = 16'b1111111110000101;
        samples[2] = 16'b1111111010100111;
        samples[3] = 16'b1111111111000000;
        samples[4] = 16'b1111110011101011;
        samples[5] = 16'b1111111101100101;
        samples[6] = 16'b0000000100000101;
        samples[7] = 16'b1111111110001000;
        samples[8] = 16'b1111110011001000;
        samples[9] = 16'b0000000000000010;
        samples[10] = 16'b0000000111101111;
        samples[11] = 16'b0000001011100011;
        samples[12] = 16'b1111110101010010;
        samples[13] = 16'b0000001000100001;
        samples[14] = 16'b0000001010011000;
        samples[15] = 16'b1111111110001110;
        samples[16] = 16'b0000001001000111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011111011;
        samples[1] = 16'b1111111110100001;
        samples[2] = 16'b1111111010111001;
        samples[3] = 16'b1111111111111011;
        samples[4] = 16'b1111110011010101;
        samples[5] = 16'b1111111110011110;
        samples[6] = 16'b0000000100000010;
        samples[7] = 16'b1111111111000110;
        samples[8] = 16'b1111110001110111;
        samples[9] = 16'b0000000100101110;
        samples[10] = 16'b0000000111011010;
        samples[11] = 16'b0000001001101100;
        samples[12] = 16'b1111110101100010;
        samples[13] = 16'b0000000001000110;
        samples[14] = 16'b0000000111100011;
        samples[15] = 16'b1111111111001100;
        samples[16] = 16'b0000001000110111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100110000;
        samples[1] = 16'b1111111111001100;
        samples[2] = 16'b1111111010001110;
        samples[3] = 16'b1111111111011111;
        samples[4] = 16'b1111110100001010;
        samples[5] = 16'b1111111110100111;
        samples[6] = 16'b0000000011011001;
        samples[7] = 16'b1111111111001100;
        samples[8] = 16'b1111110011011011;
        samples[9] = 16'b0000000011001010;
        samples[10] = 16'b0000001000000010;
        samples[11] = 16'b0000001000011110;
        samples[12] = 16'b1111111001011100;
        samples[13] = 16'b0000000100110100;
        samples[14] = 16'b0000000110110001;
        samples[15] = 16'b1111111111101100;
        samples[16] = 16'b0000001000000010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101001100;
        samples[1] = 16'b1111111110111010;
        samples[2] = 16'b1111111010001110;
        samples[3] = 16'b0000000000001110;
        samples[4] = 16'b1111110100110110;
        samples[5] = 16'b1111111110110000;
        samples[6] = 16'b0000000010101010;
        samples[7] = 16'b0000000000000010;
        samples[8] = 16'b1111110100101001;
        samples[9] = 16'b0000000010010001;
        samples[10] = 16'b0000001000100101;
        samples[11] = 16'b0000001001000111;
        samples[12] = 16'b0000000001010000;
        samples[13] = 16'b0000000101101100;
        samples[14] = 16'b0000000111101100;
        samples[15] = 16'b0000000000010100;
        samples[16] = 16'b0000000111000001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101010011;
        samples[1] = 16'b1111111101111011;
        samples[2] = 16'b1111111001111011;
        samples[3] = 16'b0000000010000010;
        samples[4] = 16'b1111110101101011;
        samples[5] = 16'b1111111110010111;
        samples[6] = 16'b0000000010000010;
        samples[7] = 16'b0000000000111101;
        samples[8] = 16'b1111110100111111;
        samples[9] = 16'b0000000110001000;
        samples[10] = 16'b0000000111110011;
        samples[11] = 16'b0000001001010111;
        samples[12] = 16'b0000000110010101;
        samples[13] = 16'b1111111101111011;
        samples[14] = 16'b0000000111000001;
        samples[15] = 16'b0000000001000011;
        samples[16] = 16'b0000000110000101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101000011;
        samples[1] = 16'b1111111101110101;
        samples[2] = 16'b1111111001000110;
        samples[3] = 16'b0000000010110111;
        samples[4] = 16'b1111110110000001;
        samples[5] = 16'b1111111101111000;
        samples[6] = 16'b0000000000011011;
        samples[7] = 16'b0000000010010100;
        samples[8] = 16'b1111111000100110;
        samples[9] = 16'b0000000100011000;
        samples[10] = 16'b0000000110000101;
        samples[11] = 16'b0000000111000001;
        samples[12] = 16'b0000000001010110;
        samples[13] = 16'b0000001011101101;
        samples[14] = 16'b0000000100010010;
        samples[15] = 16'b0000000001000000;
        samples[16] = 16'b0000000100010101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100100100;
        samples[1] = 16'b1111111101011100;
        samples[2] = 16'b1111111000111100;
        samples[3] = 16'b0000000011111100;
        samples[4] = 16'b1111110110011010;
        samples[5] = 16'b1111111101010110;
        samples[6] = 16'b1111111111010000;
        samples[7] = 16'b0000000011110010;
        samples[8] = 16'b1111111011011100;
        samples[9] = 16'b0000000011110010;
        samples[10] = 16'b0000000011110101;
        samples[11] = 16'b0000000101111001;
        samples[12] = 16'b0000000001011111;
        samples[13] = 16'b0000010010000110;
        samples[14] = 16'b0000000011000110;
        samples[15] = 16'b0000000001011100;
        samples[16] = 16'b0000000010101010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101000110;
        samples[1] = 16'b1111111100111010;
        samples[2] = 16'b1111111001111000;
        samples[3] = 16'b0000000101010000;
        samples[4] = 16'b1111110111011000;
        samples[5] = 16'b1111111101011100;
        samples[6] = 16'b0000000000001011;
        samples[7] = 16'b0000000011110101;
        samples[8] = 16'b1111111101101111;
        samples[9] = 16'b0000001001110110;
        samples[10] = 16'b0000000000101010;
        samples[11] = 16'b0000000101100110;
        samples[12] = 16'b1111111000001010;
        samples[13] = 16'b0000001000011110;
        samples[14] = 16'b0000000001011100;
        samples[15] = 16'b0000000010111101;
        samples[16] = 16'b0000000010101010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101110010;
        samples[1] = 16'b1111111101011111;
        samples[2] = 16'b1111111010111001;
        samples[3] = 16'b0000000100001011;
        samples[4] = 16'b1111111000100011;
        samples[5] = 16'b1111111110001110;
        samples[6] = 16'b0000000000110100;
        samples[7] = 16'b0000000010100100;
        samples[8] = 16'b0000000001100010;
        samples[9] = 16'b0000001000100001;
        samples[10] = 16'b1111111111101001;
        samples[11] = 16'b0000000011000011;
        samples[12] = 16'b0000000011111111;
        samples[13] = 16'b1111111111100010;
        samples[14] = 16'b1111111111011001;
        samples[15] = 16'b0000000011111100;
        samples[16] = 16'b0000000010010001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110110011;
        samples[1] = 16'b1111111110111010;
        samples[2] = 16'b1111111100000100;
        samples[3] = 16'b0000000010010001;
        samples[4] = 16'b1111111001111110;
        samples[5] = 16'b1111111111100101;
        samples[6] = 16'b0000000000011011;
        samples[7] = 16'b0000000001110010;
        samples[8] = 16'b0000000011000011;
        samples[9] = 16'b0000000110111101;
        samples[10] = 16'b0000000000001011;
        samples[11] = 16'b0000000001010011;
        samples[12] = 16'b0000000100010010;
        samples[13] = 16'b0000000001110101;
        samples[14] = 16'b1111111110010111;
        samples[15] = 16'b0000000100110111;
        samples[16] = 16'b0000000001001001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111111111011;
        samples[1] = 16'b1111111111000011;
        samples[2] = 16'b1111111100010001;
        samples[3] = 16'b0000000010111101;
        samples[4] = 16'b1111111010111100;
        samples[5] = 16'b0000000000111010;
        samples[6] = 16'b1111111111110010;
        samples[7] = 16'b0000000010011011;
        samples[8] = 16'b0000000001111011;
        samples[9] = 16'b0000000100111010;
        samples[10] = 16'b0000000010110111;
        samples[11] = 16'b0000000010101101;
        samples[12] = 16'b0000001010010010;
        samples[13] = 16'b1111111110010100;
        samples[14] = 16'b1111111111000110;
        samples[15] = 16'b0000000100111101;
        samples[16] = 16'b0000000001001101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000000111010;
        samples[1] = 16'b1111111111011100;
        samples[2] = 16'b1111111100101101;
        samples[3] = 16'b0000000010100001;
        samples[4] = 16'b1111111100001011;
        samples[5] = 16'b0000000010001000;
        samples[6] = 16'b1111111111101111;
        samples[7] = 16'b0000000001011100;
        samples[8] = 16'b0000000011111000;
        samples[9] = 16'b0000000100110001;
        samples[10] = 16'b0000000010011110;
        samples[11] = 16'b0000000001010110;
        samples[12] = 16'b0000010001100111;
        samples[13] = 16'b1111111110010001;
        samples[14] = 16'b1111111111011111;
        samples[15] = 16'b0000000101010110;
        samples[16] = 16'b0000000001010000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000001010011;
        samples[1] = 16'b1111111111011111;
        samples[2] = 16'b1111111100100001;
        samples[3] = 16'b0000000010111101;
        samples[4] = 16'b1111111100010001;
        samples[5] = 16'b0000000010110001;
        samples[6] = 16'b1111111111001001;
        samples[7] = 16'b0000000001111111;
        samples[8] = 16'b0000000011111000;
        samples[9] = 16'b0000000100101011;
        samples[10] = 16'b0000000010000010;
        samples[11] = 16'b0000000001010011;
        samples[12] = 16'b0000001010001111;
        samples[13] = 16'b0000000101001010;
        samples[14] = 16'b0000000000100100;
        samples[15] = 16'b0000000101001101;
        samples[16] = 16'b0000000000111010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000010100001;
        samples[1] = 16'b1111111111111011;
        samples[2] = 16'b1111111101011100;
        samples[3] = 16'b0000000010010100;
        samples[4] = 16'b1111111101011100;
        samples[5] = 16'b0000000011011100;
        samples[6] = 16'b1111111111001100;
        samples[7] = 16'b0000000010000010;
        samples[8] = 16'b0000000110000101;
        samples[9] = 16'b0000000011010011;
        samples[10] = 16'b0000000001110101;
        samples[11] = 16'b0000000010000101;
        samples[12] = 16'b0000000111000100;
        samples[13] = 16'b0000010111101110;
        samples[14] = 16'b0000000010000101;
        samples[15] = 16'b0000000101010000;
        samples[16] = 16'b0000000001001101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011010000;
        samples[1] = 16'b0000000000001011;
        samples[2] = 16'b1111111110000001;
        samples[3] = 16'b0000000010000101;
        samples[4] = 16'b1111111101100101;
        samples[5] = 16'b0000000011100110;
        samples[6] = 16'b0000000000001011;
        samples[7] = 16'b0000000010000101;
        samples[8] = 16'b0000000100010010;
        samples[9] = 16'b0000000100111010;
        samples[10] = 16'b0000000010110001;
        samples[11] = 16'b0000000001110010;
        samples[12] = 16'b0000001001011101;
        samples[13] = 16'b0000001011011010;
        samples[14] = 16'b0000000001101001;
        samples[15] = 16'b0000000101111001;
        samples[16] = 16'b0000000001111111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011111100;
        samples[1] = 16'b0000000000110100;
        samples[2] = 16'b1111111110001000;
        samples[3] = 16'b0000000001010011;
        samples[4] = 16'b1111111101111110;
        samples[5] = 16'b0000000100000101;
        samples[6] = 16'b0000000000101010;
        samples[7] = 16'b0000000001011100;
        samples[8] = 16'b0000000101011101;
        samples[9] = 16'b0000000010011011;
        samples[10] = 16'b0000000011100011;
        samples[11] = 16'b0000000000111101;
        samples[12] = 16'b0000001011110000;
        samples[13] = 16'b0000001100001001;
        samples[14] = 16'b0000000000001110;
        samples[15] = 16'b0000000101111111;
        samples[16] = 16'b0000000010011110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000100110001;
        samples[1] = 16'b0000000001000011;
        samples[2] = 16'b1111111110001110;
        samples[3] = 16'b0000000001011001;
        samples[4] = 16'b1111111110101101;
        samples[5] = 16'b0000000100010101;
        samples[6] = 16'b0000000000110111;
        samples[7] = 16'b0000000001011100;
        samples[8] = 16'b0000000100000010;
        samples[9] = 16'b0000000010100111;
        samples[10] = 16'b0000000100110100;
        samples[11] = 16'b0000000010110100;
        samples[12] = 16'b0000001011000100;
        samples[13] = 16'b0000001011110011;
        samples[14] = 16'b0000000010110100;
        samples[15] = 16'b0000000110100100;
        samples[16] = 16'b0000000010110100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101010000;
        samples[1] = 16'b0000000000100100;
        samples[2] = 16'b1111111110001011;
        samples[3] = 16'b0000000010011110;
        samples[4] = 16'b1111111111100101;
        samples[5] = 16'b0000000100011000;
        samples[6] = 16'b0000000001001001;
        samples[7] = 16'b0000000001001101;
        samples[8] = 16'b0000000100000010;
        samples[9] = 16'b0000000100100001;
        samples[10] = 16'b0000000100110111;
        samples[11] = 16'b0000000011000011;
        samples[12] = 16'b0000010000110101;
        samples[13] = 16'b1111101110101100;
        samples[14] = 16'b0000000001111111;
        samples[15] = 16'b0000000111101001;
        samples[16] = 16'b0000000010110100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101010110;
        samples[1] = 16'b0000000001101001;
        samples[2] = 16'b1111111111000011;
        samples[3] = 16'b0000000001100010;
        samples[4] = 16'b0000000000110000;
        samples[5] = 16'b0000000101011001;
        samples[6] = 16'b0000000001101111;
        samples[7] = 16'b1111111111101100;
        samples[8] = 16'b0000001000111010;
        samples[9] = 16'b0000000110110001;
        samples[10] = 16'b0000000010000101;
        samples[11] = 16'b1111111110100100;
        samples[12] = 16'b0000001010110100;
        samples[13] = 16'b1111110100100011;
        samples[14] = 16'b1111111111100010;
        samples[15] = 16'b0000001000100101;
        samples[16] = 16'b0000000010000010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101011101;
        samples[1] = 16'b0000000010100001;
        samples[2] = 16'b1111111111101111;
        samples[3] = 16'b0000000001011001;
        samples[4] = 16'b0000000001111000;
        samples[5] = 16'b0000000101101111;
        samples[6] = 16'b0000000001111000;
        samples[7] = 16'b1111111111011100;
        samples[8] = 16'b0000001000000101;
        samples[9] = 16'b0000000101100011;
        samples[10] = 16'b0000000011111111;
        samples[11] = 16'b1111111101110101;
        samples[12] = 16'b0000000110101011;
        samples[13] = 16'b1111111010101010;
        samples[14] = 16'b0000000000001110;
        samples[15] = 16'b0000001000111110;
        samples[16] = 16'b0000000001101111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110011011;
        samples[1] = 16'b0000000010110111;
        samples[2] = 16'b0000000001110010;
        samples[3] = 16'b0000000001100110;
        samples[4] = 16'b0000000011101001;
        samples[5] = 16'b0000000101110010;
        samples[6] = 16'b0000000011010110;
        samples[7] = 16'b1111111111111000;
        samples[8] = 16'b0000001001011101;
        samples[9] = 16'b0000000100101011;
        samples[10] = 16'b0000000101001101;
        samples[11] = 16'b1111111111111011;
        samples[12] = 16'b0000001101010100;
        samples[13] = 16'b1111110110110110;
        samples[14] = 16'b0000000010111101;
        samples[15] = 16'b0000001001110000;
        samples[16] = 16'b0000000010100111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110110111;
        samples[1] = 16'b0000000011101100;
        samples[2] = 16'b0000000011011111;
        samples[3] = 16'b0000000001100010;
        samples[4] = 16'b0000000100100111;
        samples[5] = 16'b0000000101111100;
        samples[6] = 16'b0000000101001010;
        samples[7] = 16'b1111111111111110;
        samples[8] = 16'b0000001000001111;
        samples[9] = 16'b0000000101000100;
        samples[10] = 16'b0000000111100011;
        samples[11] = 16'b0000000010001000;
        samples[12] = 16'b0000001101010111;
        samples[13] = 16'b1111110110110000;
        samples[14] = 16'b0000000101101111;
        samples[15] = 16'b0000001010011000;
        samples[16] = 16'b0000000011111100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110100001;
        samples[1] = 16'b0000000100110001;
        samples[2] = 16'b0000000100111010;
        samples[3] = 16'b0000000001111011;
        samples[4] = 16'b0000000100101110;
        samples[5] = 16'b0000000101110010;
        samples[6] = 16'b0000000101100011;
        samples[7] = 16'b0000000010000101;
        samples[8] = 16'b0000000111111001;
        samples[9] = 16'b0000000100110100;
        samples[10] = 16'b0000001000000101;
        samples[11] = 16'b0000000011000000;
        samples[12] = 16'b0000001110101000;
        samples[13] = 16'b1111111111101100;
        samples[14] = 16'b0000000110110100;
        samples[15] = 16'b0000001010101000;
        samples[16] = 16'b0000000100010010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101111111;
        samples[1] = 16'b0000000101010011;
        samples[2] = 16'b0000000111000111;
        samples[3] = 16'b0000000011001101;
        samples[4] = 16'b0000000100010101;
        samples[5] = 16'b0000000101100000;
        samples[6] = 16'b0000000110110100;
        samples[7] = 16'b0000000100111101;
        samples[8] = 16'b0000000110001111;
        samples[9] = 16'b0000001010100101;
        samples[10] = 16'b0000000110111010;
        samples[11] = 16'b0000000011101100;
        samples[12] = 16'b0000001101101010;
        samples[13] = 16'b1111111111100101;
        samples[14] = 16'b0000000110000010;
        samples[15] = 16'b0000001011110000;
        samples[16] = 16'b0000000100111010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110100100;
        samples[1] = 16'b0000000101111001;
        samples[2] = 16'b0000001000101110;
        samples[3] = 16'b0000000010100001;
        samples[4] = 16'b0000000100111010;
        samples[5] = 16'b0000000101111001;
        samples[6] = 16'b0000001000110001;
        samples[7] = 16'b0000000100001000;
        samples[8] = 16'b0000001000100001;
        samples[9] = 16'b0000001100001111;
        samples[10] = 16'b0000000101111111;
        samples[11] = 16'b0000000011110010;
        samples[12] = 16'b0000010100001001;
        samples[13] = 16'b1111111011101000;
        samples[14] = 16'b0000001000010010;
        samples[15] = 16'b0000001100110101;
        samples[16] = 16'b0000000101101001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000100110001;
        samples[1] = 16'b0000000101010000;
        samples[2] = 16'b0000001001001010;
        samples[3] = 16'b0000000100110111;
        samples[4] = 16'b0000000011100110;
        samples[5] = 16'b0000000101011101;
        samples[6] = 16'b0000001000101011;
        samples[7] = 16'b0000000110001111;
        samples[8] = 16'b0000001011101001;
        samples[9] = 16'b0000001010011110;
        samples[10] = 16'b0000000100111010;
        samples[11] = 16'b0000000011000110;
        samples[12] = 16'b0000001011010111;
        samples[13] = 16'b0000010110010110;
        samples[14] = 16'b0000000110101000;
        samples[15] = 16'b0000001100001001;
        samples[16] = 16'b0000000100110100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101010000;
        samples[1] = 16'b0000000101000111;
        samples[2] = 16'b0000001001100000;
        samples[3] = 16'b0000000101011001;
        samples[4] = 16'b0000000100000101;
        samples[5] = 16'b0000000110001111;
        samples[6] = 16'b0000000111100011;
        samples[7] = 16'b0000000111011010;
        samples[8] = 16'b0000001100100010;
        samples[9] = 16'b0000001010101110;
        samples[10] = 16'b0000000100111010;
        samples[11] = 16'b0000000011001101;
        samples[12] = 16'b0000001111011010;
        samples[13] = 16'b0000000111010110;
        samples[14] = 16'b0000000011010011;
        samples[15] = 16'b0000001011101001;
        samples[16] = 16'b0000000100100111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101111001;
        samples[1] = 16'b0000000101011101;
        samples[2] = 16'b0000001010001001;
        samples[3] = 16'b0000000100100111;
        samples[4] = 16'b0000000101000111;
        samples[5] = 16'b0000000110101110;
        samples[6] = 16'b0000000111101111;
        samples[7] = 16'b0000000110101000;
        samples[8] = 16'b0000001110111110;
        samples[9] = 16'b0000001010111011;
        samples[10] = 16'b0000000101011001;
        samples[11] = 16'b0000000010001011;
        samples[12] = 16'b0000001011100000;
        samples[13] = 16'b0000000011100110;
        samples[14] = 16'b0000000000001000;
        samples[15] = 16'b0000001011010111;
        samples[16] = 16'b0000000101010110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101000100;
        samples[1] = 16'b0000000100011011;
        samples[2] = 16'b0000001001000100;
        samples[3] = 16'b0000000110001011;
        samples[4] = 16'b0000000100000101;
        samples[5] = 16'b0000000101100000;
        samples[6] = 16'b0000000111011101;
        samples[7] = 16'b0000000111101111;
        samples[8] = 16'b0000001101000100;
        samples[9] = 16'b0000001001000100;
        samples[10] = 16'b0000000111010011;
        samples[11] = 16'b0000000010110001;
        samples[12] = 16'b0000001000111110;
        samples[13] = 16'b0000000000100100;
        samples[14] = 16'b1111111111111011;
        samples[15] = 16'b0000001001111001;
        samples[16] = 16'b0000000101001010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101100000;
        samples[1] = 16'b0000000100100111;
        samples[2] = 16'b0000001001100110;
        samples[3] = 16'b0000000101010011;
        samples[4] = 16'b0000000100101011;
        samples[5] = 16'b0000000101100110;
        samples[6] = 16'b0000000111101001;
        samples[7] = 16'b0000000111000100;
        samples[8] = 16'b0000001101111100;
        samples[9] = 16'b0000001110001100;
        samples[10] = 16'b0000000101110010;
        samples[11] = 16'b0000000000000010;
        samples[12] = 16'b0000001011000111;
        samples[13] = 16'b0000000000010111;
        samples[14] = 16'b1111111101000000;
        samples[15] = 16'b0000001001110000;
        samples[16] = 16'b0000000100110001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101101100;
        samples[1] = 16'b0000000100011011;
        samples[2] = 16'b0000001001110011;
        samples[3] = 16'b0000000100010010;
        samples[4] = 16'b0000000100100100;
        samples[5] = 16'b0000000101000100;
        samples[6] = 16'b0000000111111100;
        samples[7] = 16'b0000000110101000;
        samples[8] = 16'b0000001101011010;
        samples[9] = 16'b0000010000101000;
        samples[10] = 16'b0000000100111010;
        samples[11] = 16'b1111111111000000;
        samples[12] = 16'b0000001011111001;
        samples[13] = 16'b0000000110110111;
        samples[14] = 16'b1111111101011001;
        samples[15] = 16'b0000001001010011;
        samples[16] = 16'b0000000100010010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000100110001;
        samples[1] = 16'b0000000011010011;
        samples[2] = 16'b0000001000110001;
        samples[3] = 16'b0000000100101011;
        samples[4] = 16'b0000000011101001;
        samples[5] = 16'b0000000011100011;
        samples[6] = 16'b0000000110110111;
        samples[7] = 16'b0000000111100011;
        samples[8] = 16'b0000010011000001;
        samples[9] = 16'b0000001001100000;
        samples[10] = 16'b0000000001110010;
        samples[11] = 16'b1111111101100010;
        samples[12] = 16'b0000001100011100;
        samples[13] = 16'b0000000101000000;
        samples[14] = 16'b1111111101011001;
        samples[15] = 16'b0000000111001101;
        samples[16] = 16'b0000000010010001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000100100100;
        samples[1] = 16'b0000000011011001;
        samples[2] = 16'b0000001000100101;
        samples[3] = 16'b0000000011000011;
        samples[4] = 16'b0000000011100110;
        samples[5] = 16'b0000000011010110;
        samples[6] = 16'b0000000101111001;
        samples[7] = 16'b0000000110110100;
        samples[8] = 16'b0000010100100010;
        samples[9] = 16'b0000001011011101;
        samples[10] = 16'b1111111111100101;
        samples[11] = 16'b1111111001001001;
        samples[12] = 16'b0000001011110011;
        samples[13] = 16'b0000001011010000;
        samples[14] = 16'b1111110110110110;
        samples[15] = 16'b0000000110011000;
        samples[16] = 16'b0000000000110111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101010000;
        samples[1] = 16'b0000000011101100;
        samples[2] = 16'b0000000111011101;
        samples[3] = 16'b0000000001011100;
        samples[4] = 16'b0000000100010101;
        samples[5] = 16'b0000000010101010;
        samples[6] = 16'b0000000100100100;
        samples[7] = 16'b0000000110001111;
        samples[8] = 16'b0000010111000101;
        samples[9] = 16'b0000000111100011;
        samples[10] = 16'b1111111101110101;
        samples[11] = 16'b1111111001101011;
        samples[12] = 16'b0000001111111101;
        samples[13] = 16'b0000001101110110;
        samples[14] = 16'b1111111000110011;
        samples[15] = 16'b0000000101000100;
        samples[16] = 16'b1111111111011100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101111001;
        samples[1] = 16'b0000000011011001;
        samples[2] = 16'b0000000110001011;
        samples[3] = 16'b1111111111110010;
        samples[4] = 16'b0000000100101011;
        samples[5] = 16'b0000000001011111;
        samples[6] = 16'b0000000011111000;
        samples[7] = 16'b0000000101000100;
        samples[8] = 16'b0000010101101101;
        samples[9] = 16'b0000000100101110;
        samples[10] = 16'b1111111110100100;
        samples[11] = 16'b1111111010111100;
        samples[12] = 16'b0000001100011100;
        samples[13] = 16'b0000010001001000;
        samples[14] = 16'b1111111001001001;
        samples[15] = 16'b0000000011101111;
        samples[16] = 16'b1111111110001110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101010000;
        samples[1] = 16'b0000000011101001;
        samples[2] = 16'b0000000100101011;
        samples[3] = 16'b1111111110110000;
        samples[4] = 16'b0000000100000010;
        samples[5] = 16'b0000000000100001;
        samples[6] = 16'b0000000010101101;
        samples[7] = 16'b0000000100111101;
        samples[8] = 16'b0000010001110110;
        samples[9] = 16'b0000000011111100;
        samples[10] = 16'b0000000000001110;
        samples[11] = 16'b1111111000111111;
        samples[12] = 16'b0000010010011100;
        samples[13] = 16'b0000001001001101;
        samples[14] = 16'b1111110110010100;
        samples[15] = 16'b0000000001111000;
        samples[16] = 16'b1111111101000000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000100100100;
        samples[1] = 16'b0000000011001010;
        samples[2] = 16'b0000000011000011;
        samples[3] = 16'b1111111111000011;
        samples[4] = 16'b0000000011111111;
        samples[5] = 16'b1111111111010011;
        samples[6] = 16'b0000000001010000;
        samples[7] = 16'b0000000101011001;
        samples[8] = 16'b0000010100000110;
        samples[9] = 16'b0000000000011011;
        samples[10] = 16'b1111111101101111;
        samples[11] = 16'b1111110111100101;
        samples[12] = 16'b0000010110110101;
        samples[13] = 16'b0000001110101000;
        samples[14] = 16'b1111110110111111;
        samples[15] = 16'b1111111111101001;
        samples[16] = 16'b1111111011101000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011010110;
        samples[1] = 16'b0000000001010110;
        samples[2] = 16'b0000000001011111;
        samples[3] = 16'b0000000000000010;
        samples[4] = 16'b0000000011001010;
        samples[5] = 16'b1111111101100101;
        samples[6] = 16'b0000000000110000;
        samples[7] = 16'b0000000100110100;
        samples[8] = 16'b0000010110000110;
        samples[9] = 16'b1111111110110011;
        samples[10] = 16'b1111111001100101;
        samples[11] = 16'b1111110111100010;
        samples[12] = 16'b0000010010111011;
        samples[13] = 16'b0000000000001011;
        samples[14] = 16'b1111110101110100;
        samples[15] = 16'b1111111101011001;
        samples[16] = 16'b1111111010111001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000001010011;
        samples[1] = 16'b0000000000001011;
        samples[2] = 16'b0000000000010001;
        samples[3] = 16'b0000000001000000;
        samples[4] = 16'b0000000001110101;
        samples[5] = 16'b1111111100001011;
        samples[6] = 16'b0000000000011110;
        samples[7] = 16'b0000000100011011;
        samples[8] = 16'b0000010110010011;
        samples[9] = 16'b1111111110010001;
        samples[10] = 16'b1111110111110001;
        samples[11] = 16'b1111110101110100;
        samples[12] = 16'b0000010010110101;
        samples[13] = 16'b1111111111011111;
        samples[14] = 16'b1111110011111010;
        samples[15] = 16'b1111111011110101;
        samples[16] = 16'b1111111010001010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110110111;
        samples[1] = 16'b1111111111100010;
        samples[2] = 16'b1111111111100010;
        samples[3] = 16'b0000000010001000;
        samples[4] = 16'b1111111111111110;
        samples[5] = 16'b1111111011000000;
        samples[6] = 16'b1111111111010011;
        samples[7] = 16'b0000000101101111;
        samples[8] = 16'b0000010101011011;
        samples[9] = 16'b1111111101001100;
        samples[10] = 16'b1111110101101110;
        samples[11] = 16'b1111110010111100;
        samples[12] = 16'b0000000111100110;
        samples[13] = 16'b0000000001101001;
        samples[14] = 16'b1111101111100100;
        samples[15] = 16'b1111111010101101;
        samples[16] = 16'b1111111000111001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101011001;
        samples[1] = 16'b1111111110110111;
        samples[2] = 16'b1111111111000110;
        samples[3] = 16'b0000000010011011;
        samples[4] = 16'b1111111110011110;
        samples[5] = 16'b1111111010011101;
        samples[6] = 16'b1111111111011111;
        samples[7] = 16'b0000000101011001;
        samples[8] = 16'b0000010000111000;
        samples[9] = 16'b1111111101010011;
        samples[10] = 16'b1111110110010100;
        samples[11] = 16'b1111110011010010;
        samples[12] = 16'b0000000100001000;
        samples[13] = 16'b0000001100000011;
        samples[14] = 16'b1111110000011100;
        samples[15] = 16'b1111111010010111;
        samples[16] = 16'b1111111001010010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100010111;
        samples[1] = 16'b1111111110011010;
        samples[2] = 16'b1111111110100111;
        samples[3] = 16'b0000000010001110;
        samples[4] = 16'b1111111101000000;
        samples[5] = 16'b1111111010100000;
        samples[6] = 16'b0000000000011011;
        samples[7] = 16'b0000000011011100;
        samples[8] = 16'b0000001100101000;
        samples[9] = 16'b1111111101100101;
        samples[10] = 16'b1111111001100010;
        samples[11] = 16'b1111110010101111;
        samples[12] = 16'b1111111111101001;
        samples[13] = 16'b0000000100100100;
        samples[14] = 16'b1111110000110101;
        samples[15] = 16'b1111111010110011;
        samples[16] = 16'b1111111010010100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100001110;
        samples[1] = 16'b1111111110001011;
        samples[2] = 16'b1111111111001100;
        samples[3] = 16'b0000000010011110;
        samples[4] = 16'b1111111100101101;
        samples[5] = 16'b1111111011111110;
        samples[6] = 16'b0000000000010111;
        samples[7] = 16'b0000000010110111;
        samples[8] = 16'b0000001100001001;
        samples[9] = 16'b1111111000010100;
        samples[10] = 16'b1111111100001011;
        samples[11] = 16'b1111110011111010;
        samples[12] = 16'b0000001100111000;
        samples[13] = 16'b1111110101101000;
        samples[14] = 16'b1111110011101110;
        samples[15] = 16'b1111111001101110;
        samples[16] = 16'b1111111011101011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100100111;
        samples[1] = 16'b1111111110110111;
        samples[2] = 16'b1111111111000000;
        samples[3] = 16'b0000000001000110;
        samples[4] = 16'b1111111100001110;
        samples[5] = 16'b1111111101001111;
        samples[6] = 16'b0000000000001011;
        samples[7] = 16'b0000000001101111;
        samples[8] = 16'b0000000111010011;
        samples[9] = 16'b1111110111000010;
        samples[10] = 16'b1111111110010100;
        samples[11] = 16'b1111110110101101;
        samples[12] = 16'b0000001101110011;
        samples[13] = 16'b1111111000000001;
        samples[14] = 16'b1111110111111000;
        samples[15] = 16'b1111111001010101;
        samples[16] = 16'b1111111101011001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100000100;
        samples[1] = 16'b1111111111000000;
        samples[2] = 16'b1111111110101010;
        samples[3] = 16'b0000000001111011;
        samples[4] = 16'b1111111011011001;
        samples[5] = 16'b1111111101110101;
        samples[6] = 16'b0000000000010111;
        samples[7] = 16'b0000000001111111;
        samples[8] = 16'b0000001001010011;
        samples[9] = 16'b1111110010101001;
        samples[10] = 16'b1111111110011010;
        samples[11] = 16'b1111111000000111;
        samples[12] = 16'b0000001010011011;
        samples[13] = 16'b1111110000110101;
        samples[14] = 16'b1111110110110011;
        samples[15] = 16'b1111111000100110;
        samples[16] = 16'b1111111110011010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011111011;
        samples[1] = 16'b1111111111111011;
        samples[2] = 16'b1111111111100010;
        samples[3] = 16'b0000000001100010;
        samples[4] = 16'b1111111010111001;
        samples[5] = 16'b1111111111101001;
        samples[6] = 16'b0000000000111010;
        samples[7] = 16'b0000000001010011;
        samples[8] = 16'b0000000110100001;
        samples[9] = 16'b1111110100111001;
        samples[10] = 16'b1111111111100101;
        samples[11] = 16'b1111110111101011;
        samples[12] = 16'b0000000111100011;
        samples[13] = 16'b1111110010000000;
        samples[14] = 16'b1111110101011110;
        samples[15] = 16'b1111111001001100;
        samples[16] = 16'b0000000000000010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011100101;
        samples[1] = 16'b0000000000011011;
        samples[2] = 16'b1111111111011111;
        samples[3] = 16'b0000000001011111;
        samples[4] = 16'b1111111010000100;
        samples[5] = 16'b0000000000010001;
        samples[6] = 16'b0000000001010110;
        samples[7] = 16'b0000000001010000;
        samples[8] = 16'b0000000010001110;
        samples[9] = 16'b1111110101011110;
        samples[10] = 16'b0000000001101100;
        samples[11] = 16'b1111111001011000;
        samples[12] = 16'b0000000011111111;
        samples[13] = 16'b0000000001011100;
        samples[14] = 16'b1111110111100010;
        samples[15] = 16'b1111111001111000;
        samples[16] = 16'b0000000000111101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011110101;
        samples[1] = 16'b0000000000011110;
        samples[2] = 16'b1111111111001100;
        samples[3] = 16'b0000000001110010;
        samples[4] = 16'b1111111001111110;
        samples[5] = 16'b0000000000110100;
        samples[6] = 16'b0000000001011001;
        samples[7] = 16'b0000000001000000;
        samples[8] = 16'b1111111110001000;
        samples[9] = 16'b1111110101110100;
        samples[10] = 16'b0000000100111101;
        samples[11] = 16'b1111111011000000;
        samples[12] = 16'b0000001001000001;
        samples[13] = 16'b1111110101001100;
        samples[14] = 16'b1111110111000010;
        samples[15] = 16'b1111111010110011;
        samples[16] = 16'b0000000001111000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100000001;
        samples[1] = 16'b0000000000011011;
        samples[2] = 16'b1111111111011001;
        samples[3] = 16'b0000000010000010;
        samples[4] = 16'b1111111010110000;
        samples[5] = 16'b0000000001011001;
        samples[6] = 16'b0000000000110111;
        samples[7] = 16'b0000000000110000;
        samples[8] = 16'b0000000000001011;
        samples[9] = 16'b1111110111010101;
        samples[10] = 16'b0000000010110001;
        samples[11] = 16'b1111111001011111;
        samples[12] = 16'b1111111111110101;
        samples[13] = 16'b1111111011010101;
        samples[14] = 16'b1111111000001010;
        samples[15] = 16'b1111111011101000;
        samples[16] = 16'b0000000001100010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100001011;
        samples[1] = 16'b0000000000100100;
        samples[2] = 16'b1111111110110111;
        samples[3] = 16'b0000000001111011;
        samples[4] = 16'b1111111011000110;
        samples[5] = 16'b0000000001100010;
        samples[6] = 16'b0000000000001110;
        samples[7] = 16'b0000000000100100;
        samples[8] = 16'b1111111101110101;
        samples[9] = 16'b1111111000010100;
        samples[10] = 16'b0000000011101100;
        samples[11] = 16'b1111111001001100;
        samples[12] = 16'b0000000000010100;
        samples[13] = 16'b0000001000011000;
        samples[14] = 16'b1111111010011101;
        samples[15] = 16'b1111111100100100;
        samples[16] = 16'b0000000001000011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101011100;
        samples[1] = 16'b0000000000010111;
        samples[2] = 16'b1111111111000011;
        samples[3] = 16'b0000000001010000;
        samples[4] = 16'b1111111101001111;
        samples[5] = 16'b0000000001111111;
        samples[6] = 16'b1111111111110101;
        samples[7] = 16'b1111111110111101;
        samples[8] = 16'b1111111101111011;
        samples[9] = 16'b1111111011010101;
        samples[10] = 16'b0000000011010011;
        samples[11] = 16'b1111111001001001;
        samples[12] = 16'b1111111100010100;
        samples[13] = 16'b1111111110010100;
        samples[14] = 16'b1111111010011010;
        samples[15] = 16'b1111111110001011;
        samples[16] = 16'b0000000000111101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110101101;
        samples[1] = 16'b0000000000001110;
        samples[2] = 16'b1111111111011001;
        samples[3] = 16'b0000000000101010;
        samples[4] = 16'b1111111111010011;
        samples[5] = 16'b0000000010100111;
        samples[6] = 16'b1111111111101100;
        samples[7] = 16'b1111111101010011;
        samples[8] = 16'b1111111110101101;
        samples[9] = 16'b1111111111000000;
        samples[10] = 16'b0000000001101111;
        samples[11] = 16'b1111111000111001;
        samples[12] = 16'b1111110110100000;
        samples[13] = 16'b0000000001111111;
        samples[14] = 16'b1111111100001011;
        samples[15] = 16'b1111111111001100;
        samples[16] = 16'b0000000000111010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110000001;
        samples[1] = 16'b1111111111111000;
        samples[2] = 16'b1111111111000011;
        samples[3] = 16'b0000000001100110;
        samples[4] = 16'b1111111111010000;
        samples[5] = 16'b0000000010101010;
        samples[6] = 16'b1111111110101101;
        samples[7] = 16'b1111111101110101;
        samples[8] = 16'b1111111011001111;
        samples[9] = 16'b0000000000010001;
        samples[10] = 16'b0000000010111010;
        samples[11] = 16'b1111111000001101;
        samples[12] = 16'b1111111010110011;
        samples[13] = 16'b0000000100000101;
        samples[14] = 16'b1111111010111001;
        samples[15] = 16'b1111111111011001;
        samples[16] = 16'b0000000000010100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110000001;
        samples[1] = 16'b0000000000011110;
        samples[2] = 16'b0000000000010111;
        samples[3] = 16'b0000000000011110;
        samples[4] = 16'b0000000000100001;
        samples[5] = 16'b0000000010111010;
        samples[6] = 16'b1111111111000000;
        samples[7] = 16'b1111111100111010;
        samples[8] = 16'b1111111100100001;
        samples[9] = 16'b1111111101111000;
        samples[10] = 16'b0000000011101001;
        samples[11] = 16'b1111110111010101;
        samples[12] = 16'b0000000111001010;
        samples[13] = 16'b1111101110111100;
        samples[14] = 16'b1111111000001101;
        samples[15] = 16'b1111111111010110;
        samples[16] = 16'b0000000000000101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110000001;
        samples[1] = 16'b0000000000001110;
        samples[2] = 16'b0000000001000000;
        samples[3] = 16'b0000000000101101;
        samples[4] = 16'b0000000000110100;
        samples[5] = 16'b0000000010100111;
        samples[6] = 16'b0000000000000010;
        samples[7] = 16'b1111111100100001;
        samples[8] = 16'b1111111011000110;
        samples[9] = 16'b1111111111000011;
        samples[10] = 16'b0000000011110010;
        samples[11] = 16'b1111111001011100;
        samples[12] = 16'b0000000100100111;
        samples[13] = 16'b1111111001100010;
        samples[14] = 16'b1111111011001100;
        samples[15] = 16'b0000000000000010;
        samples[16] = 16'b0000000000010100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100100100;
        samples[1] = 16'b1111111111110101;
        samples[2] = 16'b0000000001011111;
        samples[3] = 16'b0000000001111011;
        samples[4] = 16'b1111111111111000;
        samples[5] = 16'b0000000001011100;
        samples[6] = 16'b0000000000100111;
        samples[7] = 16'b1111111101101111;
        samples[8] = 16'b1111111000100000;
        samples[9] = 16'b1111111110001011;
        samples[10] = 16'b0000000011111100;
        samples[11] = 16'b1111111100010111;
        samples[12] = 16'b0000001001000100;
        samples[13] = 16'b1111111000001101;
        samples[14] = 16'b1111111101011111;
        samples[15] = 16'b1111111111101111;
        samples[16] = 16'b1111111111101001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011101110;
        samples[1] = 16'b0000000001000110;
        samples[2] = 16'b0000000011000110;
        samples[3] = 16'b1111111111110010;
        samples[4] = 16'b1111111111111011;
        samples[5] = 16'b0000000001010110;
        samples[6] = 16'b0000000001001001;
        samples[7] = 16'b1111111101001100;
        samples[8] = 16'b1111111010100011;
        samples[9] = 16'b1111111101111000;
        samples[10] = 16'b0000000001111000;
        samples[11] = 16'b1111111001100101;
        samples[12] = 16'b0000001010001111;
        samples[13] = 16'b1111111010001010;
        samples[14] = 16'b1111111100001011;
        samples[15] = 16'b1111111111101001;
        samples[16] = 16'b1111111110010100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011000011;
        samples[1] = 16'b0000000001100010;
        samples[2] = 16'b0000000011110101;
        samples[3] = 16'b1111111111000000;
        samples[4] = 16'b1111111111100010;
        samples[5] = 16'b0000000001011100;
        samples[6] = 16'b0000000001100010;
        samples[7] = 16'b1111111100111010;
        samples[8] = 16'b1111110110010111;
        samples[9] = 16'b0000000000000101;
        samples[10] = 16'b0000000011110010;
        samples[11] = 16'b1111111001001100;
        samples[12] = 16'b1111111010010111;
        samples[13] = 16'b0000001011111001;
        samples[14] = 16'b1111111010010001;
        samples[15] = 16'b1111111111100010;
        samples[16] = 16'b1111111110110111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111010110000;
        samples[1] = 16'b0000000001000000;
        samples[2] = 16'b0000000011011111;
        samples[3] = 16'b1111111111000011;
        samples[4] = 16'b1111111111000000;
        samples[5] = 16'b0000000001000110;
        samples[6] = 16'b0000000001100010;
        samples[7] = 16'b1111111100100111;
        samples[8] = 16'b1111110101110100;
        samples[9] = 16'b1111111000110110;
        samples[10] = 16'b0000000110111010;
        samples[11] = 16'b1111111011010010;
        samples[12] = 16'b1111111101011001;
        samples[13] = 16'b1111111101000011;
        samples[14] = 16'b1111111101110101;
        samples[15] = 16'b1111111101001111;
        samples[16] = 16'b1111111111000011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111001101000;
        samples[1] = 16'b0000000001000000;
        samples[2] = 16'b0000000100001000;
        samples[3] = 16'b1111111111100010;
        samples[4] = 16'b1111111110110111;
        samples[5] = 16'b0000000001010011;
        samples[6] = 16'b0000000001011100;
        samples[7] = 16'b1111111100101101;
        samples[8] = 16'b1111111010000001;
        samples[9] = 16'b1111111001000110;
        samples[10] = 16'b0000000011111000;
        samples[11] = 16'b1111111000110000;
        samples[12] = 16'b1111111010010100;
        samples[13] = 16'b1111111011001111;
        samples[14] = 16'b1111111100010001;
        samples[15] = 16'b1111111100100001;
        samples[16] = 16'b1111111110110111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111001001111;
        samples[1] = 16'b0000000001011001;
        samples[2] = 16'b0000000101011001;
        samples[3] = 16'b1111111110111010;
        samples[4] = 16'b1111111111010000;
        samples[5] = 16'b0000000001101111;
        samples[6] = 16'b0000000001011111;
        samples[7] = 16'b1111111100010100;
        samples[8] = 16'b1111111100000100;
        samples[9] = 16'b1111111010101010;
        samples[10] = 16'b0000000001111011;
        samples[11] = 16'b1111111000010111;
        samples[12] = 16'b1111110110010000;
        samples[13] = 16'b1111111101100101;
        samples[14] = 16'b1111111011000000;
        samples[15] = 16'b1111111100010111;
        samples[16] = 16'b1111111110110011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111000110011;
        samples[1] = 16'b0000000001110101;
        samples[2] = 16'b0000000110000101;
        samples[3] = 16'b1111111101111110;
        samples[4] = 16'b1111111110100111;
        samples[5] = 16'b0000000001111000;
        samples[6] = 16'b0000000010001000;
        samples[7] = 16'b1111111100000100;
        samples[8] = 16'b1111111010101101;
        samples[9] = 16'b1111111011111011;
        samples[10] = 16'b0000000001011100;
        samples[11] = 16'b1111111001010010;
        samples[12] = 16'b1111110001110001;
        samples[13] = 16'b0000001000000101;
        samples[14] = 16'b1111111110000001;
        samples[15] = 16'b1111111100111010;
        samples[16] = 16'b1111111110110011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111101110;
        samples[1] = 16'b0000000010011000;
        samples[2] = 16'b0000000110011011;
        samples[3] = 16'b1111111110000001;
        samples[4] = 16'b1111111101111110;
        samples[5] = 16'b0000000001111111;
        samples[6] = 16'b0000000010000010;
        samples[7] = 16'b1111111100100001;
        samples[8] = 16'b1111111011011001;
        samples[9] = 16'b1111111011000000;
        samples[10] = 16'b1111111110001110;
        samples[11] = 16'b1111111000000100;
        samples[12] = 16'b1111111000100110;
        samples[13] = 16'b0000000100100001;
        samples[14] = 16'b1111111111000000;
        samples[15] = 16'b1111111100111101;
        samples[16] = 16'b1111111101101111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111110100;
        samples[1] = 16'b0000000011000011;
        samples[2] = 16'b0000000111010000;
        samples[3] = 16'b1111111100010001;
        samples[4] = 16'b1111111101010011;
        samples[5] = 16'b0000000010100001;
        samples[6] = 16'b0000000010101101;
        samples[7] = 16'b1111111011101110;
        samples[8] = 16'b1111111000011101;
        samples[9] = 16'b1111111010110000;
        samples[10] = 16'b0000000000001110;
        samples[11] = 16'b1111111000111001;
        samples[12] = 16'b0000000000000010;
        samples[13] = 16'b0000000010100100;
        samples[14] = 16'b1111111111000000;
        samples[15] = 16'b1111111101101111;
        samples[16] = 16'b1111111101110101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111111011;
        samples[1] = 16'b0000000010011110;
        samples[2] = 16'b0000000110010101;
        samples[3] = 16'b1111111101001100;
        samples[4] = 16'b1111111100001110;
        samples[5] = 16'b0000000010010001;
        samples[6] = 16'b0000000010101101;
        samples[7] = 16'b1111111100110000;
        samples[8] = 16'b1111110110110110;
        samples[9] = 16'b1111110110110110;
        samples[10] = 16'b0000000011000011;
        samples[11] = 16'b1111111011110101;
        samples[12] = 16'b1111111111101111;
        samples[13] = 16'b1111111111011100;
        samples[14] = 16'b1111111111111000;
        samples[15] = 16'b1111111101100010;
        samples[16] = 16'b1111111110011110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111000000001;
        samples[1] = 16'b0000000010000010;
        samples[2] = 16'b0000000101001101;
        samples[3] = 16'b1111111110010001;
        samples[4] = 16'b1111111011010101;
        samples[5] = 16'b0000000001111111;
        samples[6] = 16'b0000000010011000;
        samples[7] = 16'b1111111101101100;
        samples[8] = 16'b1111111000000100;
        samples[9] = 16'b1111110111000010;
        samples[10] = 16'b0000000010011000;
        samples[11] = 16'b1111111010110011;
        samples[12] = 16'b0000000010011000;
        samples[13] = 16'b1111110101101011;
        samples[14] = 16'b1111111101111011;
        samples[15] = 16'b1111111101011111;
        samples[16] = 16'b1111111111000011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111111110;
        samples[1] = 16'b0000000010010001;
        samples[2] = 16'b0000000100110100;
        samples[3] = 16'b1111111110100001;
        samples[4] = 16'b1111111011011001;
        samples[5] = 16'b0000000010100111;
        samples[6] = 16'b0000000010000101;
        samples[7] = 16'b1111111101011100;
        samples[8] = 16'b1111111111111011;
        samples[9] = 16'b1111111011011111;
        samples[10] = 16'b1111111011001001;
        samples[11] = 16'b1111110110100011;
        samples[12] = 16'b1111111100010001;
        samples[13] = 16'b1111111001000011;
        samples[14] = 16'b1111111001010010;
        samples[15] = 16'b1111111101111000;
        samples[16] = 16'b1111111110110111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111001100101;
        samples[1] = 16'b0000000010100111;
        samples[2] = 16'b0000000100110001;
        samples[3] = 16'b1111111100100100;
        samples[4] = 16'b1111111100001110;
        samples[5] = 16'b0000000011100011;
        samples[6] = 16'b0000000010100100;
        samples[7] = 16'b1111111011001001;
        samples[8] = 16'b0000000011010000;
        samples[9] = 16'b1111111011000011;
        samples[10] = 16'b1111111010110110;
        samples[11] = 16'b1111110111001111;
        samples[12] = 16'b1111111100011101;
        samples[13] = 16'b1111110011000101;
        samples[14] = 16'b1111111010100011;
        samples[15] = 16'b1111111110100100;
        samples[16] = 16'b1111111111100101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111001110101;
        samples[1] = 16'b0000000010000101;
        samples[2] = 16'b0000000011101100;
        samples[3] = 16'b1111111101000110;
        samples[4] = 16'b1111111011011111;
        samples[5] = 16'b0000000011011111;
        samples[6] = 16'b0000000010010100;
        samples[7] = 16'b1111111011010010;
        samples[8] = 16'b0000000000001011;
        samples[9] = 16'b1111111001011000;
        samples[10] = 16'b1111111100001011;
        samples[11] = 16'b1111111010010001;
        samples[12] = 16'b1111111111100010;
        samples[13] = 16'b1111110001011000;
        samples[14] = 16'b1111111101101111;
        samples[15] = 16'b1111111110011110;
        samples[16] = 16'b1111111111101001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111010000100;
        samples[1] = 16'b0000000010110001;
        samples[2] = 16'b0000000011000000;
        samples[3] = 16'b1111111011001100;
        samples[4] = 16'b1111111010110011;
        samples[5] = 16'b0000000011110101;
        samples[6] = 16'b0000000001101111;
        samples[7] = 16'b1111111010101010;
        samples[8] = 16'b1111111100010111;
        samples[9] = 16'b1111111001001111;
        samples[10] = 16'b1111111101111110;
        samples[11] = 16'b1111111001001001;
        samples[12] = 16'b0000000001101100;
        samples[13] = 16'b1111110000010110;
        samples[14] = 16'b1111111101010110;
        samples[15] = 16'b1111111110110000;
        samples[16] = 16'b1111111110111101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111001111110;
        samples[1] = 16'b0000000010101010;
        samples[2] = 16'b0000000001101001;
        samples[3] = 16'b1111111011001100;
        samples[4] = 16'b1111111001011000;
        samples[5] = 16'b0000000011001010;
        samples[6] = 16'b0000000001001101;
        samples[7] = 16'b1111111011110010;
        samples[8] = 16'b1111110101101011;
        samples[9] = 16'b1111111100010100;
        samples[10] = 16'b1111111111111110;
        samples[11] = 16'b1111111010010111;
        samples[12] = 16'b1111111100100111;
        samples[13] = 16'b1111101111011000;
        samples[14] = 16'b1111111100111010;
        samples[15] = 16'b1111111111101001;
        samples[16] = 16'b1111111110111101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111010000001;
        samples[1] = 16'b0000000010000010;
        samples[2] = 16'b0000000000001110;
        samples[3] = 16'b1111111100110110;
        samples[4] = 16'b1111111000101101;
        samples[5] = 16'b0000000001111000;
        samples[6] = 16'b0000000001111111;
        samples[7] = 16'b1111111100011101;
        samples[8] = 16'b1111110111111110;
        samples[9] = 16'b1111111101110101;
        samples[10] = 16'b1111111110010111;
        samples[11] = 16'b1111111100000100;
        samples[12] = 16'b1111110101011011;
        samples[13] = 16'b0000000011101111;
        samples[14] = 16'b1111111010100111;
        samples[15] = 16'b0000000000000101;
        samples[16] = 16'b1111111111011001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111010011010;
        samples[1] = 16'b0000000010100100;
        samples[2] = 16'b0000000000011110;
        samples[3] = 16'b1111111010111001;
        samples[4] = 16'b1111111000111111;
        samples[5] = 16'b0000000001110010;
        samples[6] = 16'b0000000010110001;
        samples[7] = 16'b1111111010110110;
        samples[8] = 16'b1111111010011101;
        samples[9] = 16'b0000000000100111;
        samples[10] = 16'b1111111100001110;
        samples[11] = 16'b1111111000111111;
        samples[12] = 16'b1111111100001000;
        samples[13] = 16'b1111111111011100;
        samples[14] = 16'b1111111001101000;
        samples[15] = 16'b0000000000010100;
        samples[16] = 16'b1111111111011111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111001001001;
        samples[1] = 16'b0000000010110100;
        samples[2] = 16'b0000000000100100;
        samples[3] = 16'b1111111011011001;
        samples[4] = 16'b1111111000010001;
        samples[5] = 16'b0000000001011111;
        samples[6] = 16'b0000000010000010;
        samples[7] = 16'b1111111100001000;
        samples[8] = 16'b0000000000100001;
        samples[9] = 16'b1111111110001110;
        samples[10] = 16'b1111111000100011;
        samples[11] = 16'b1111110110011010;
        samples[12] = 16'b1111110000110010;
        samples[13] = 16'b0000001010001100;
        samples[14] = 16'b1111110100110000;
        samples[15] = 16'b1111111111100010;
        samples[16] = 16'b1111111110010100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111010010111;
        samples[1] = 16'b0000000011101100;
        samples[2] = 16'b0000000001010000;
        samples[3] = 16'b1111111001110001;
        samples[4] = 16'b1111111001011111;
        samples[5] = 16'b0000000010010001;
        samples[6] = 16'b0000000010001011;
        samples[7] = 16'b1111111011001100;
        samples[8] = 16'b1111111111000110;
        samples[9] = 16'b1111111011100010;
        samples[10] = 16'b1111111100110000;
        samples[11] = 16'b1111110111101011;
        samples[12] = 16'b1111111010001010;
        samples[13] = 16'b0000001000010101;
        samples[14] = 16'b1111110101110001;
        samples[15] = 16'b1111111111000011;
        samples[16] = 16'b1111111110110111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111001011100;
        samples[1] = 16'b0000000010110001;
        samples[2] = 16'b0000000001000110;
        samples[3] = 16'b1111111100001110;
        samples[4] = 16'b1111111000011010;
        samples[5] = 16'b0000000001001101;
        samples[6] = 16'b0000000010000010;
        samples[7] = 16'b1111111101111000;
        samples[8] = 16'b1111111010000001;
        samples[9] = 16'b1111111011000110;
        samples[10] = 16'b1111111111011001;
        samples[11] = 16'b1111111001000110;
        samples[12] = 16'b0000000100111101;
        samples[13] = 16'b0000000000001011;
        samples[14] = 16'b1111111001111011;
        samples[15] = 16'b1111111110011010;
        samples[16] = 16'b1111111110100111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111001111110;
        samples[1] = 16'b0000000010011110;
        samples[2] = 16'b0000000001000110;
        samples[3] = 16'b1111111100100111;
        samples[4] = 16'b1111111000101101;
        samples[5] = 16'b0000000000101010;
        samples[6] = 16'b0000000001111000;
        samples[7] = 16'b1111111110110111;
        samples[8] = 16'b1111110011100001;
        samples[9] = 16'b1111111101000110;
        samples[10] = 16'b0000000011110101;
        samples[11] = 16'b1111111010101010;
        samples[12] = 16'b1111111011001001;
        samples[13] = 16'b1111111010101010;
        samples[14] = 16'b1111111010000001;
        samples[15] = 16'b1111111111101111;
        samples[16] = 16'b1111111110101010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111010111100;
        samples[1] = 16'b0000000010111101;
        samples[2] = 16'b0000000001101111;
        samples[3] = 16'b1111111101000011;
        samples[4] = 16'b1111111010000100;
        samples[5] = 16'b0000000000101101;
        samples[6] = 16'b0000000010000010;
        samples[7] = 16'b1111111111110101;
        samples[8] = 16'b1111110111010010;
        samples[9] = 16'b1111111101111110;
        samples[10] = 16'b0000000011100011;
        samples[11] = 16'b1111111011111110;
        samples[12] = 16'b1111111100010001;
        samples[13] = 16'b1111111000111100;
        samples[14] = 16'b1111111001100101;
        samples[15] = 16'b0000000000111010;
        samples[16] = 16'b1111111110100100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111100000001;
        samples[1] = 16'b0000000011000000;
        samples[2] = 16'b0000000010010001;
        samples[3] = 16'b1111111101101100;
        samples[4] = 16'b1111111011010101;
        samples[5] = 16'b0000000000000101;
        samples[6] = 16'b0000000010110100;
        samples[7] = 16'b0000000000101010;
        samples[8] = 16'b1111111000001101;
        samples[9] = 16'b0000000000010001;
        samples[10] = 16'b0000000001110101;
        samples[11] = 16'b1111111100001110;
        samples[12] = 16'b0000000101111111;
        samples[13] = 16'b1111110000011100;
        samples[14] = 16'b1111111011101011;
        samples[15] = 16'b0000000001100010;
        samples[16] = 16'b1111111110100111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101011001;
        samples[1] = 16'b0000000100000101;
        samples[2] = 16'b0000000011101001;
        samples[3] = 16'b1111111100110000;
        samples[4] = 16'b1111111100110011;
        samples[5] = 16'b0000000000101010;
        samples[6] = 16'b0000000011111100;
        samples[7] = 16'b0000000000010001;
        samples[8] = 16'b1111111001111011;
        samples[9] = 16'b1111111111000011;
        samples[10] = 16'b0000000100011011;
        samples[11] = 16'b1111111011001001;
        samples[12] = 16'b1111111101101000;
        samples[13] = 16'b1111111000111111;
        samples[14] = 16'b1111110111101011;
        samples[15] = 16'b0000000010001011;
        samples[16] = 16'b1111111111111000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110000001;
        samples[1] = 16'b0000000100011011;
        samples[2] = 16'b0000000100100001;
        samples[3] = 16'b1111111101100010;
        samples[4] = 16'b1111111101111110;
        samples[5] = 16'b0000000000110100;
        samples[6] = 16'b0000000100100111;
        samples[7] = 16'b0000000001000011;
        samples[8] = 16'b1111111010100111;
        samples[9] = 16'b0000000100100111;
        samples[10] = 16'b0000000001010011;
        samples[11] = 16'b1111111100100100;
        samples[12] = 16'b1111111101000000;
        samples[13] = 16'b0000001010111011;
        samples[14] = 16'b1111111001011000;
        samples[15] = 16'b0000000010001110;
        samples[16] = 16'b0000000000010111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110011110;
        samples[1] = 16'b0000000011001101;
        samples[2] = 16'b0000000100100001;
        samples[3] = 16'b0000000000101010;
        samples[4] = 16'b1111111110011110;
        samples[5] = 16'b1111111111101111;
        samples[6] = 16'b0000000100111010;
        samples[7] = 16'b0000000011101100;
        samples[8] = 16'b1111111001010101;
        samples[9] = 16'b0000000100000101;
        samples[10] = 16'b0000000000111101;
        samples[11] = 16'b0000000000011011;
        samples[12] = 16'b0000001011110000;
        samples[13] = 16'b1111111001010101;
        samples[14] = 16'b1111111100101010;
        samples[15] = 16'b0000000001011001;
        samples[16] = 16'b0000000000111010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110100111;
        samples[1] = 16'b0000000011000011;
        samples[2] = 16'b0000000101010110;
        samples[3] = 16'b0000000001000110;
        samples[4] = 16'b1111111110100100;
        samples[5] = 16'b1111111111101111;
        samples[6] = 16'b0000000101101100;
        samples[7] = 16'b0000000100000101;
        samples[8] = 16'b1111110111000010;
        samples[9] = 16'b0000000101000000;
        samples[10] = 16'b0000000010110100;
        samples[11] = 16'b1111111111101111;
        samples[12] = 16'b1111111010111100;
        samples[13] = 16'b0000001110101110;
        samples[14] = 16'b1111111001111011;
        samples[15] = 16'b0000000001101111;
        samples[16] = 16'b0000000001011001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110011010;
        samples[1] = 16'b0000000010100001;
        samples[2] = 16'b0000000101010000;
        samples[3] = 16'b0000000010100100;
        samples[4] = 16'b1111111110100100;
        samples[5] = 16'b1111111111011001;
        samples[6] = 16'b0000000101001101;
        samples[7] = 16'b0000000101100011;
        samples[8] = 16'b1111110111111000;
        samples[9] = 16'b0000000001010011;
        samples[10] = 16'b0000000010100111;
        samples[11] = 16'b0000000001001101;
        samples[12] = 16'b0000000000110111;
        samples[13] = 16'b1111111011110101;
        samples[14] = 16'b1111111010011010;
        samples[15] = 16'b0000000001100010;
        samples[16] = 16'b0000000000101101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000000000010;
        samples[1] = 16'b0000000010011110;
        samples[2] = 16'b0000000110011110;
        samples[3] = 16'b0000000010011000;
        samples[4] = 16'b0000000000001011;
        samples[5] = 16'b0000000000001000;
        samples[6] = 16'b0000000101111111;
        samples[7] = 16'b0000000101000100;
        samples[8] = 16'b1111111110011010;
        samples[9] = 16'b0000000000101101;
        samples[10] = 16'b1111111111101001;
        samples[11] = 16'b0000000010100111;
        samples[12] = 16'b0000001111101101;
        samples[13] = 16'b1111101111111101;
        samples[14] = 16'b1111111101111000;
        samples[15] = 16'b0000000010001110;
        samples[16] = 16'b0000000000010100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000000110000;
        samples[1] = 16'b0000000010100111;
        samples[2] = 16'b0000000110110100;
        samples[3] = 16'b0000000001100010;
        samples[4] = 16'b0000000000100100;
        samples[5] = 16'b0000000000010001;
        samples[6] = 16'b0000000110110100;
        samples[7] = 16'b0000000100001011;
        samples[8] = 16'b1111111100110011;
        samples[9] = 16'b1111111111011100;
        samples[10] = 16'b0000000010100111;
        samples[11] = 16'b0000000011110010;
        samples[12] = 16'b0000000111100011;
        samples[13] = 16'b1111110100100110;
        samples[14] = 16'b1111111101000011;
        samples[15] = 16'b0000000011000110;
        samples[16] = 16'b0000000000101101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000001000110;
        samples[1] = 16'b0000000011010011;
        samples[2] = 16'b0000000110101011;
        samples[3] = 16'b0000000000110100;
        samples[4] = 16'b0000000000010100;
        samples[5] = 16'b0000000000000010;
        samples[6] = 16'b0000000110010010;
        samples[7] = 16'b0000000101001101;
        samples[8] = 16'b1111111001111000;
        samples[9] = 16'b1111111111101100;
        samples[10] = 16'b0000000101001101;
        samples[11] = 16'b0000000011111000;
        samples[12] = 16'b0000001111000100;
        samples[13] = 16'b1111111011101110;
        samples[14] = 16'b1111111011011100;
        samples[15] = 16'b0000000011011100;
        samples[16] = 16'b0000000000010001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000000111101;
        samples[1] = 16'b0000000010001011;
        samples[2] = 16'b0000000101000100;
        samples[3] = 16'b0000000010100001;
        samples[4] = 16'b1111111111011100;
        samples[5] = 16'b1111111110010001;
        samples[6] = 16'b0000000101001010;
        samples[7] = 16'b0000000111111100;
        samples[8] = 16'b1111110111110100;
        samples[9] = 16'b0000000010011000;
        samples[10] = 16'b0000000100001011;
        samples[11] = 16'b0000000100100001;
        samples[12] = 16'b0000001110000000;
        samples[13] = 16'b0000000011011111;
        samples[14] = 16'b1111111011000000;
        samples[15] = 16'b0000000011001101;
        samples[16] = 16'b1111111111101001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000001100010;
        samples[1] = 16'b0000000000101010;
        samples[2] = 16'b0000000011000011;
        samples[3] = 16'b0000000011100110;
        samples[4] = 16'b1111111110111101;
        samples[5] = 16'b1111111101001001;
        samples[6] = 16'b0000000100110111;
        samples[7] = 16'b0000000111111111;
        samples[8] = 16'b1111110101110100;
        samples[9] = 16'b0000000010011110;
        samples[10] = 16'b0000000110001011;
        samples[11] = 16'b0000000101111001;
        samples[12] = 16'b0000000010111101;
        samples[13] = 16'b0000001110001111;
        samples[14] = 16'b1111111100101101;
        samples[15] = 16'b0000000100000101;
        samples[16] = 16'b0000000000001011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011001010;
        samples[1] = 16'b0000000000101010;
        samples[2] = 16'b0000000010011110;
        samples[3] = 16'b0000000010011000;
        samples[4] = 16'b0000000000001000;
        samples[5] = 16'b1111111110000001;
        samples[6] = 16'b0000000100101011;
        samples[7] = 16'b0000000101111100;
        samples[8] = 16'b1111111000110011;
        samples[9] = 16'b0000000011110010;
        samples[10] = 16'b0000000110111101;
        samples[11] = 16'b0000000100001011;
        samples[12] = 16'b0000000100100100;
        samples[13] = 16'b0000011110101001;
        samples[14] = 16'b1111111011111011;
        samples[15] = 16'b0000000100100001;
        samples[16] = 16'b0000000000010111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011111000;
        samples[1] = 16'b1111111111101111;
        samples[2] = 16'b0000000000100100;
        samples[3] = 16'b0000000011010110;
        samples[4] = 16'b0000000000000010;
        samples[5] = 16'b1111111110100001;
        samples[6] = 16'b0000000010000101;
        samples[7] = 16'b0000000111000100;
        samples[8] = 16'b1111111001011000;
        samples[9] = 16'b0000000011111000;
        samples[10] = 16'b0000000101101100;
        samples[11] = 16'b0000000101100000;
        samples[12] = 16'b0000000111100000;
        samples[13] = 16'b0000010001000100;
        samples[14] = 16'b1111111110110111;
        samples[15] = 16'b0000000011111100;
        samples[16] = 16'b1111111111101100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000100111010;
        samples[1] = 16'b0000000000101010;
        samples[2] = 16'b0000000000100111;
        samples[3] = 16'b0000000001111011;
        samples[4] = 16'b0000000000110000;
        samples[5] = 16'b0000000000000101;
        samples[6] = 16'b0000000010010001;
        samples[7] = 16'b0000000101001010;
        samples[8] = 16'b1111111010010100;
        samples[9] = 16'b0000000110001000;
        samples[10] = 16'b0000000111110110;
        samples[11] = 16'b0000000011111100;
        samples[12] = 16'b0000001101100000;
        samples[13] = 16'b0000001011010100;
        samples[14] = 16'b1111111001101110;
        samples[15] = 16'b0000000101000111;
        samples[16] = 16'b0000000000110000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101010000;
        samples[1] = 16'b0000000001011111;
        samples[2] = 16'b0000000000001011;
        samples[3] = 16'b0000000001011001;
        samples[4] = 16'b0000000001010110;
        samples[5] = 16'b0000000000100111;
        samples[6] = 16'b0000000010010100;
        samples[7] = 16'b0000000100001000;
        samples[8] = 16'b1111111100110110;
        samples[9] = 16'b0000000000100001;
        samples[10] = 16'b0000001001111111;
        samples[11] = 16'b0000000011011100;
        samples[12] = 16'b0000010010010011;
        samples[13] = 16'b1111111111101001;
        samples[14] = 16'b1111111001101110;
        samples[15] = 16'b0000000100011011;
        samples[16] = 16'b0000000001000011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101000100;
        samples[1] = 16'b0000000001011111;
        samples[2] = 16'b1111111111011001;
        samples[3] = 16'b0000000010011000;
        samples[4] = 16'b0000000001000110;
        samples[5] = 16'b0000000000100111;
        samples[6] = 16'b0000000001100010;
        samples[7] = 16'b0000000101000000;
        samples[8] = 16'b1111110111101011;
        samples[9] = 16'b0000000011010011;
        samples[10] = 16'b0000001011001101;
        samples[11] = 16'b0000000011111100;
        samples[12] = 16'b0000010000100010;
        samples[13] = 16'b1111111110111010;
        samples[14] = 16'b1111111011111011;
        samples[15] = 16'b0000000100100001;
        samples[16] = 16'b0000000001001001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101110110;
        samples[1] = 16'b0000000010011000;
        samples[2] = 16'b1111111111111110;
        samples[3] = 16'b0000000001010011;
        samples[4] = 16'b0000000010111101;
        samples[5] = 16'b0000000001101111;
        samples[6] = 16'b0000000001100110;
        samples[7] = 16'b0000000011001101;
        samples[8] = 16'b1111111111010000;
        samples[9] = 16'b0000001001010000;
        samples[10] = 16'b0000000100000010;
        samples[11] = 16'b0000000000101010;
        samples[12] = 16'b0000000001011100;
        samples[13] = 16'b0000000010000101;
        samples[14] = 16'b1111111010111001;
        samples[15] = 16'b0000000101110110;
        samples[16] = 16'b0000000001000110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110011110;
        samples[1] = 16'b0000000011000011;
        samples[2] = 16'b0000000000010100;
        samples[3] = 16'b0000000000000010;
        samples[4] = 16'b0000000100010010;
        samples[5] = 16'b0000000010101010;
        samples[6] = 16'b0000000001110010;
        samples[7] = 16'b0000000001001101;
        samples[8] = 16'b0000000010011011;
        samples[9] = 16'b0000001000101011;
        samples[10] = 16'b0000000010100111;
        samples[11] = 16'b1111111111000011;
        samples[12] = 16'b1111111101101100;
        samples[13] = 16'b0000000011101100;
        samples[14] = 16'b1111111011111110;
        samples[15] = 16'b0000000110000010;
        samples[16] = 16'b0000000000101101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110011000;
        samples[1] = 16'b0000000011000000;
        samples[2] = 16'b0000000000010100;
        samples[3] = 16'b0000000000010001;
        samples[4] = 16'b0000000101010011;
        samples[5] = 16'b0000000011010000;
        samples[6] = 16'b0000000000101101;
        samples[7] = 16'b0000000000110000;
        samples[8] = 16'b0000000101111100;
        samples[9] = 16'b0000000110000010;
        samples[10] = 16'b0000000001010000;
        samples[11] = 16'b1111111101011111;
        samples[12] = 16'b1111111000100110;
        samples[13] = 16'b0000010111111010;
        samples[14] = 16'b1111111011111110;
        samples[15] = 16'b0000000101101001;
        samples[16] = 16'b0000000000010001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000111000100;
        samples[1] = 16'b0000000011010011;
        samples[2] = 16'b0000000000101101;
        samples[3] = 16'b1111111111001001;
        samples[4] = 16'b0000000110110111;
        samples[5] = 16'b0000000011111100;
        samples[6] = 16'b0000000000010111;
        samples[7] = 16'b1111111111000110;
        samples[8] = 16'b0000000110001011;
        samples[9] = 16'b0000000111011010;
        samples[10] = 16'b0000000001011100;
        samples[11] = 16'b1111111101111011;
        samples[12] = 16'b0000000001101111;
        samples[13] = 16'b0000010010101100;
        samples[14] = 16'b1111111010010111;
        samples[15] = 16'b0000000110000010;
        samples[16] = 16'b0000000000000010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110111101;
        samples[1] = 16'b0000000010101101;
        samples[2] = 16'b0000000000010100;
        samples[3] = 16'b1111111110110011;
        samples[4] = 16'b0000000111000001;
        samples[5] = 16'b0000000011011111;
        samples[6] = 16'b1111111111111110;
        samples[7] = 16'b1111111110011110;
        samples[8] = 16'b0000000010101010;
        samples[9] = 16'b0000000001110010;
        samples[10] = 16'b0000000110011110;
        samples[11] = 16'b0000000000111010;
        samples[12] = 16'b0000010010100010;
        samples[13] = 16'b0000000001010011;
        samples[14] = 16'b1111111110011010;
        samples[15] = 16'b0000000101100011;
        samples[16] = 16'b1111111111101111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101101100;
        samples[1] = 16'b0000000001111011;
        samples[2] = 16'b1111111111101100;
        samples[3] = 16'b0000000000000010;
        samples[4] = 16'b0000000110011000;
        samples[5] = 16'b0000000010110100;
        samples[6] = 16'b1111111110100100;
        samples[7] = 16'b1111111111100101;
        samples[8] = 16'b1111111110000101;
        samples[9] = 16'b0000000000100001;
        samples[10] = 16'b0000001000101011;
        samples[11] = 16'b0000000000000010;
        samples[12] = 16'b0000011000110010;
        samples[13] = 16'b0000000110101011;
        samples[14] = 16'b1111111110010111;
        samples[15] = 16'b0000000100101110;
        samples[16] = 16'b1111111111000011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000100111010;
        samples[1] = 16'b0000000001011100;
        samples[2] = 16'b1111111110110111;
        samples[3] = 16'b0000000000100111;
        samples[4] = 16'b0000000101111100;
        samples[5] = 16'b0000000010011110;
        samples[6] = 16'b1111111100101101;
        samples[7] = 16'b0000000000110000;
        samples[8] = 16'b1111111010001010;
        samples[9] = 16'b0000000011111000;
        samples[10] = 16'b0000001000001111;
        samples[11] = 16'b1111111111000000;
        samples[12] = 16'b0000010100010011;
        samples[13] = 16'b1111111000101010;
        samples[14] = 16'b1111111110010100;
        samples[15] = 16'b0000000100001110;
        samples[16] = 16'b1111111110011010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101111001;
        samples[1] = 16'b0000000001001001;
        samples[2] = 16'b1111111110111010;
        samples[3] = 16'b1111111111000000;
        samples[4] = 16'b0000000110101110;
        samples[5] = 16'b0000000010011110;
        samples[6] = 16'b1111111100101010;
        samples[7] = 16'b1111111111000110;
        samples[8] = 16'b1111111101001100;
        samples[9] = 16'b0000000101101001;
        samples[10] = 16'b0000000100011000;
        samples[11] = 16'b1111111110001011;
        samples[12] = 16'b0000001011000001;
        samples[13] = 16'b0000001110100010;
        samples[14] = 16'b1111111110110011;
        samples[15] = 16'b0000000100010010;
        samples[16] = 16'b1111111110001011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101110010;
        samples[1] = 16'b0000000001111111;
        samples[2] = 16'b1111111111110010;
        samples[3] = 16'b1111111110100111;
        samples[4] = 16'b0000001000101011;
        samples[5] = 16'b0000000010111010;
        samples[6] = 16'b1111111100110000;
        samples[7] = 16'b1111111101110010;
        samples[8] = 16'b0000001001001101;
        samples[9] = 16'b0000000001111011;
        samples[10] = 16'b1111111111010000;
        samples[11] = 16'b1111111011001001;
        samples[12] = 16'b0000000000111101;
        samples[13] = 16'b0000010110001101;
        samples[14] = 16'b1111111011011100;
        samples[15] = 16'b0000000011101001;
        samples[16] = 16'b1111111101100010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101110010;
        samples[1] = 16'b0000000100011011;
        samples[2] = 16'b0000000000000101;
        samples[3] = 16'b1111111101110010;
        samples[4] = 16'b0000001010000010;
        samples[5] = 16'b0000000011100110;
        samples[6] = 16'b1111111011100101;
        samples[7] = 16'b1111111111000000;
        samples[8] = 16'b0000001100010010;
        samples[9] = 16'b0000000001101001;
        samples[10] = 16'b1111111100100100;
        samples[11] = 16'b1111111001001001;
        samples[12] = 16'b1111111001101011;
        samples[13] = 16'b0000011100110000;
        samples[14] = 16'b1111110111001100;
        samples[15] = 16'b0000000011000011;
        samples[16] = 16'b1111111100010001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000111001101;
        samples[1] = 16'b0000000110001111;
        samples[2] = 16'b0000000001000000;
        samples[3] = 16'b1111111010110011;
        samples[4] = 16'b0000001011101101;
        samples[5] = 16'b0000000100011011;
        samples[6] = 16'b1111111011111000;
        samples[7] = 16'b1111111101010110;
        samples[8] = 16'b0000001010001100;
        samples[9] = 16'b0000000100011011;
        samples[10] = 16'b1111111101000011;
        samples[11] = 16'b1111111000010111;
        samples[12] = 16'b0000000101100110;
        samples[13] = 16'b0000001001110000;
        samples[14] = 16'b1111110110100110;
        samples[15] = 16'b0000000100000010;
        samples[16] = 16'b1111111100001011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110101110;
        samples[1] = 16'b0000000111000111;
        samples[2] = 16'b0000000001010110;
        samples[3] = 16'b1111111011011111;
        samples[4] = 16'b0000001100101110;
        samples[5] = 16'b0000000101000111;
        samples[6] = 16'b1111111100010100;
        samples[7] = 16'b1111111100101010;
        samples[8] = 16'b0000001101000001;
        samples[9] = 16'b0000000101010011;
        samples[10] = 16'b1111111100001000;
        samples[11] = 16'b1111110110010000;
        samples[12] = 16'b0000001111100100;
        samples[13] = 16'b1111101101010001;
        samples[14] = 16'b1111111000100011;
        samples[15] = 16'b0000000100000101;
        samples[16] = 16'b1111111100000100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000001000011110;
        samples[1] = 16'b0000001000110001;
        samples[2] = 16'b0000000001010011;
        samples[3] = 16'b1111111000101010;
        samples[4] = 16'b0000001110001111;
        samples[5] = 16'b0000000110101110;
        samples[6] = 16'b1111111011111000;
        samples[7] = 16'b1111111010011101;
        samples[8] = 16'b0000000110001011;
        samples[9] = 16'b0000000111011101;
        samples[10] = 16'b0000000001101111;
        samples[11] = 16'b1111110110010000;
        samples[12] = 16'b0000001000000101;
        samples[13] = 16'b1111110111001100;
        samples[14] = 16'b1111111011101000;
        samples[15] = 16'b0000000100011110;
        samples[16] = 16'b1111111100100111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000001001000111;
        samples[1] = 16'b0000001001010111;
        samples[2] = 16'b0000000000110111;
        samples[3] = 16'b1111110110110110;
        samples[4] = 16'b0000001110101110;
        samples[5] = 16'b0000000110110100;
        samples[6] = 16'b1111111010110011;
        samples[7] = 16'b1111111001111011;
        samples[8] = 16'b0000000110000010;
        samples[9] = 16'b0000001000001111;
        samples[10] = 16'b0000000000101101;
        samples[11] = 16'b1111110111000010;
        samples[12] = 16'b0000000111110110;
        samples[13] = 16'b1111111111010110;
        samples[14] = 16'b1111111110100001;
        samples[15] = 16'b0000000011111100;
        samples[16] = 16'b1111111011100010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000001001001010;
        samples[1] = 16'b0000001010101110;
        samples[2] = 16'b0000000001000011;
        samples[3] = 16'b1111110101001001;
        samples[4] = 16'b0000001111111001;
        samples[5] = 16'b0000000110110111;
        samples[6] = 16'b1111111011000110;
        samples[7] = 16'b1111111000010100;
        samples[8] = 16'b0000001011010111;
        samples[9] = 16'b0000000011010011;
        samples[10] = 16'b0000000000111010;
        samples[11] = 16'b1111110111110100;
        samples[12] = 16'b0000000111101100;
        samples[13] = 16'b1111111110010100;
        samples[14] = 16'b1111111111001001;
        samples[15] = 16'b0000000011001010;
        samples[16] = 16'b1111111011001100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000001001010011;
        samples[1] = 16'b0000001011100011;
        samples[2] = 16'b0000000000111101;
        samples[3] = 16'b1111110100111001;
        samples[4] = 16'b0000010001000001;
        samples[5] = 16'b0000000111000111;
        samples[6] = 16'b1111111011000011;
        samples[7] = 16'b1111110111101110;
        samples[8] = 16'b0000010011010111;
        samples[9] = 16'b0000000001000000;
        samples[10] = 16'b1111111100100001;
        samples[11] = 16'b1111110111010101;
        samples[12] = 16'b0000000001100010;
        samples[13] = 16'b0000100000010001;
        samples[14] = 16'b1111111110101101;
        samples[15] = 16'b0000000010101010;
        samples[16] = 16'b1111111010100000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000001000011110;
        samples[1] = 16'b0000001010110100;
        samples[2] = 16'b0000000000000010;
        samples[3] = 16'b1111110101110100;
        samples[4] = 16'b0000001111110011;
        samples[5] = 16'b0000000110001011;
        samples[6] = 16'b1111111010100111;
        samples[7] = 16'b1111111000110000;
        samples[8] = 16'b0000010001110110;
        samples[9] = 16'b1111111110000101;
        samples[10] = 16'b1111111101011100;
        samples[11] = 16'b1111111001011100;
        samples[12] = 16'b0000001100101011;
        samples[13] = 16'b0000000100100001;
        samples[14] = 16'b1111111101001001;
        samples[15] = 16'b0000000010001000;
        samples[16] = 16'b1111111010000001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000001000101110;
        samples[1] = 16'b0000001010010010;
        samples[2] = 16'b0000000000000010;
        samples[3] = 16'b1111110101110001;
        samples[4] = 16'b0000001111111001;
        samples[5] = 16'b0000000110001011;
        samples[6] = 16'b1111111011010010;
        samples[7] = 16'b1111110111100010;
        samples[8] = 16'b0000010011011110;
        samples[9] = 16'b0000000001111000;
        samples[10] = 16'b1111111011011001;
        samples[11] = 16'b1111111000010001;
        samples[12] = 16'b0000011110000001;
        samples[13] = 16'b1111110000101100;
        samples[14] = 16'b1111111010001110;
        samples[15] = 16'b0000000010111101;
        samples[16] = 16'b1111111010010111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000111100110;
        samples[1] = 16'b0000001001000001;
        samples[2] = 16'b1111111111100101;
        samples[3] = 16'b1111110110100000;
        samples[4] = 16'b0000001101101101;
        samples[5] = 16'b0000000101010110;
        samples[6] = 16'b1111111011101011;
        samples[7] = 16'b1111111000000111;
        samples[8] = 16'b0000001101110110;
        samples[9] = 16'b0000000001110010;
        samples[10] = 16'b1111111101011111;
        samples[11] = 16'b1111110111011000;
        samples[12] = 16'b0000010001101101;
        samples[13] = 16'b0000001010110001;
        samples[14] = 16'b1111111010101101;
        samples[15] = 16'b0000000011000000;
        samples[16] = 16'b1111111010111100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110110111;
        samples[1] = 16'b0000000111101111;
        samples[2] = 16'b1111111110100111;
        samples[3] = 16'b1111110111001111;
        samples[4] = 16'b0000001011101101;
        samples[5] = 16'b0000000100000010;
        samples[6] = 16'b1111111011011111;
        samples[7] = 16'b1111111001010101;
        samples[8] = 16'b0000001010011011;
        samples[9] = 16'b0000000010100100;
        samples[10] = 16'b1111111110110111;
        samples[11] = 16'b1111110110011010;
        samples[12] = 16'b0000000111111100;
        samples[13] = 16'b0000010000011111;
        samples[14] = 16'b1111111000110011;
        samples[15] = 16'b0000000011000011;
        samples[16] = 16'b1111111010011101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110110001;
        samples[1] = 16'b0000000111111100;
        samples[2] = 16'b1111111111010110;
        samples[3] = 16'b1111110101101000;
        samples[4] = 16'b0000001011101101;
        samples[5] = 16'b0000000100000101;
        samples[6] = 16'b1111111100010111;
        samples[7] = 16'b1111110111100010;
        samples[8] = 16'b0000010000111011;
        samples[9] = 16'b0000000011011100;
        samples[10] = 16'b1111111010100000;
        samples[11] = 16'b1111110100100011;
        samples[12] = 16'b0000001111000001;
        samples[13] = 16'b1111110111010101;
        samples[14] = 16'b1111111000111001;
        samples[15] = 16'b0000000011010110;
        samples[16] = 16'b1111111001101000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110100100;
        samples[1] = 16'b0000000111111111;
        samples[2] = 16'b0000000000001011;
        samples[3] = 16'b1111110101010101;
        samples[4] = 16'b0000001011100011;
        samples[5] = 16'b0000000100100111;
        samples[6] = 16'b1111111101010011;
        samples[7] = 16'b1111110110101101;
        samples[8] = 16'b0000010101111101;
        samples[9] = 16'b0000000011011100;
        samples[10] = 16'b1111111000010001;
        samples[11] = 16'b1111110011100100;
        samples[12] = 16'b0000001111100100;
        samples[13] = 16'b1111111011010101;
        samples[14] = 16'b1111110111100101;
        samples[15] = 16'b0000000011101001;
        samples[16] = 16'b1111111001010101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101100011;
        samples[1] = 16'b0000001000011000;
        samples[2] = 16'b0000000000001000;
        samples[3] = 16'b1111110111010010;
        samples[4] = 16'b0000001010100010;
        samples[5] = 16'b0000000101000000;
        samples[6] = 16'b1111111100110110;
        samples[7] = 16'b1111111001000011;
        samples[8] = 16'b0000011001011011;
        samples[9] = 16'b0000000101001010;
        samples[10] = 16'b1111110101001100;
        samples[11] = 16'b1111110000111001;
        samples[12] = 16'b0000001100111110;
        samples[13] = 16'b0000000001011111;
        samples[14] = 16'b1111110001111101;
        samples[15] = 16'b0000000011001101;
        samples[16] = 16'b1111111000110000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101101001;
        samples[1] = 16'b0000001001100000;
        samples[2] = 16'b0000000000111101;
        samples[3] = 16'b1111110110001010;
        samples[4] = 16'b0000001010110111;
        samples[5] = 16'b0000000110000010;
        samples[6] = 16'b1111111100111101;
        samples[7] = 16'b1111111000100110;
        samples[8] = 16'b0000011110011010;
        samples[9] = 16'b0000000110000101;
        samples[10] = 16'b1111110000100000;
        samples[11] = 16'b1111101110011111;
        samples[12] = 16'b0000100000010111;
        samples[13] = 16'b1111110010001101;
        samples[14] = 16'b1111110000001101;
        samples[15] = 16'b0000000010101101;
        samples[16] = 16'b1111111000100011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101100110;
        samples[1] = 16'b0000001000110100;
        samples[2] = 16'b0000000001000011;
        samples[3] = 16'b1111110111101000;
        samples[4] = 16'b0000001001101001;
        samples[5] = 16'b0000000101110010;
        samples[6] = 16'b1111111101111011;
        samples[7] = 16'b1111111001111000;
        samples[8] = 16'b0000011100000100;
        samples[9] = 16'b0000000100100100;
        samples[10] = 16'b1111110001100001;
        samples[11] = 16'b1111110001101110;
        samples[12] = 16'b0000001110111000;
        samples[13] = 16'b0000010110011111;
        samples[14] = 16'b1111110100110110;
        samples[15] = 16'b0000000010011000;
        samples[16] = 16'b1111111001101000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101000000;
        samples[1] = 16'b0000000111101111;
        samples[2] = 16'b0000000000010111;
        samples[3] = 16'b1111111001101011;
        samples[4] = 16'b0000000111110011;
        samples[5] = 16'b0000000100011110;
        samples[6] = 16'b1111111101110101;
        samples[7] = 16'b1111111100110011;
        samples[8] = 16'b0000010100111111;
        samples[9] = 16'b0000000001110010;
        samples[10] = 16'b1111110101000101;
        samples[11] = 16'b1111110110000100;
        samples[12] = 16'b0000001010110100;
        samples[13] = 16'b0000011111101000;
        samples[14] = 16'b1111110111111011;
        samples[15] = 16'b0000000001100010;
        samples[16] = 16'b1111111001110001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000100010101;
        samples[1] = 16'b0000000111101100;
        samples[2] = 16'b0000000000010100;
        samples[3] = 16'b1111111001000011;
        samples[4] = 16'b0000000111000100;
        samples[5] = 16'b0000000011111000;
        samples[6] = 16'b1111111100111010;
        samples[7] = 16'b1111111101100101;
        samples[8] = 16'b0000010111011011;
        samples[9] = 16'b1111111110110111;
        samples[10] = 16'b1111110011001011;
        samples[11] = 16'b1111110101010010;
        samples[12] = 16'b0000001000110100;
        samples[13] = 16'b0000010111101110;
        samples[14] = 16'b1111111010000111;
        samples[15] = 16'b0000000001000000;
        samples[16] = 16'b1111110111111011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011111000;
        samples[1] = 16'b0000000110101011;
        samples[2] = 16'b1111111111010110;
        samples[3] = 16'b1111111001100010;
        samples[4] = 16'b0000000110011000;
        samples[5] = 16'b0000000011010011;
        samples[6] = 16'b1111111011101110;
        samples[7] = 16'b1111111110000001;
        samples[8] = 16'b0000010100010011;
        samples[9] = 16'b1111111010100011;
        samples[10] = 16'b1111110110111100;
        samples[11] = 16'b1111110101110001;
        samples[12] = 16'b0000001110001001;
        samples[13] = 16'b0000001110010101;
        samples[14] = 16'b1111111000110000;
        samples[15] = 16'b1111111111111110;
        samples[16] = 16'b1111110110111001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000100111101;
        samples[1] = 16'b0000000110011110;
        samples[2] = 16'b1111111110100111;
        samples[3] = 16'b1111111001000011;
        samples[4] = 16'b0000000111111001;
        samples[5] = 16'b0000000100001000;
        samples[6] = 16'b1111111011010010;
        samples[7] = 16'b1111111011101110;
        samples[8] = 16'b0000010010001100;
        samples[9] = 16'b1111111011000000;
        samples[10] = 16'b1111111001100010;
        samples[11] = 16'b1111110100101001;
        samples[12] = 16'b0000011001110111;
        samples[13] = 16'b0000000111111111;
        samples[14] = 16'b1111110101011110;
        samples[15] = 16'b1111111111011100;
        samples[16] = 16'b1111110110100000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011111111;
        samples[1] = 16'b0000000100111101;
        samples[2] = 16'b1111111101101100;
        samples[3] = 16'b1111111100000001;
        samples[4] = 16'b0000001000000101;
        samples[5] = 16'b0000000011111100;
        samples[6] = 16'b1111111010000100;
        samples[7] = 16'b1111111100011101;
        samples[8] = 16'b0000010100000011;
        samples[9] = 16'b1111111111001100;
        samples[10] = 16'b1111110110000100;
        samples[11] = 16'b1111110010000000;
        samples[12] = 16'b0000011100111001;
        samples[13] = 16'b0000010001001110;
        samples[14] = 16'b1111101111000010;
        samples[15] = 16'b1111111110111101;
        samples[16] = 16'b1111110101101110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000100110111;
        samples[1] = 16'b0000000100011000;
        samples[2] = 16'b1111111101011001;
        samples[3] = 16'b1111111011010101;
        samples[4] = 16'b0000001001110110;
        samples[5] = 16'b0000000011111000;
        samples[6] = 16'b1111111001010010;
        samples[7] = 16'b1111111010111001;
        samples[8] = 16'b0000010010000110;
        samples[9] = 16'b1111111101110101;
        samples[10] = 16'b1111111000010100;
        samples[11] = 16'b1111110010110010;
        samples[12] = 16'b0000011101011011;
        samples[13] = 16'b0000010010010110;
        samples[14] = 16'b1111101101100100;
        samples[15] = 16'b1111111110001000;
        samples[16] = 16'b1111110101111011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000100110100;
        samples[1] = 16'b0000000011010011;
        samples[2] = 16'b1111111100110011;
        samples[3] = 16'b1111111101000011;
        samples[4] = 16'b0000001010101110;
        samples[5] = 16'b0000000011000110;
        samples[6] = 16'b1111111001000011;
        samples[7] = 16'b1111111011001001;
        samples[8] = 16'b0000001111000001;
        samples[9] = 16'b0000000000001011;
        samples[10] = 16'b1111111001011000;
        samples[11] = 16'b1111110011010010;
        samples[12] = 16'b0000101000000010;
        samples[13] = 16'b0000000111110110;
        samples[14] = 16'b1111101011111010;
        samples[15] = 16'b1111111101101111;
        samples[16] = 16'b1111110110100000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011011111;
        samples[1] = 16'b0000000001010011;
        samples[2] = 16'b1111111100110110;
        samples[3] = 16'b1111111110111101;
        samples[4] = 16'b0000001010000101;
        samples[5] = 16'b0000000001000000;
        samples[6] = 16'b1111111000110000;
        samples[7] = 16'b1111111100110011;
        samples[8] = 16'b0000001110111011;
        samples[9] = 16'b0000000000000010;
        samples[10] = 16'b1111110110110011;
        samples[11] = 16'b1111110011101000;
        samples[12] = 16'b0000011000100011;
        samples[13] = 16'b0000000001010110;
        samples[14] = 16'b1111101110010011;
        samples[15] = 16'b1111111100110000;
        samples[16] = 16'b1111110110101001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011010110;
        samples[1] = 16'b0000000000001110;
        samples[2] = 16'b1111111100111101;
        samples[3] = 16'b1111111111011001;
        samples[4] = 16'b0000001010011000;
        samples[5] = 16'b1111111111011111;
        samples[6] = 16'b1111111000111100;
        samples[7] = 16'b1111111101001111;
        samples[8] = 16'b0000010000000011;
        samples[9] = 16'b1111111111100101;
        samples[10] = 16'b1111110101010101;
        samples[11] = 16'b1111110101001111;
        samples[12] = 16'b0000011010011101;
        samples[13] = 16'b0000000110010010;
        samples[14] = 16'b1111110001101110;
        samples[15] = 16'b1111111100000100;
        samples[16] = 16'b1111110110111001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011101001;
        samples[1] = 16'b1111111110011110;
        samples[2] = 16'b1111111101001100;
        samples[3] = 16'b1111111110011010;
        samples[4] = 16'b0000001001110011;
        samples[5] = 16'b1111111101111110;
        samples[6] = 16'b1111111001110001;
        samples[7] = 16'b1111111100010001;
        samples[8] = 16'b0000010000011111;
        samples[9] = 16'b1111111010100000;
        samples[10] = 16'b1111110110001101;
        samples[11] = 16'b1111110111101110;
        samples[12] = 16'b0000001010001111;
        samples[13] = 16'b0000001101101010;
        samples[14] = 16'b1111110101011011;
        samples[15] = 16'b1111111010100011;
        samples[16] = 16'b1111110111000110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000010001110;
        samples[1] = 16'b1111111101001111;
        samples[2] = 16'b1111111101011100;
        samples[3] = 16'b0000000000000101;
        samples[4] = 16'b0000000111110011;
        samples[5] = 16'b1111111100111010;
        samples[6] = 16'b1111111010100111;
        samples[7] = 16'b1111111101110010;
        samples[8] = 16'b0000010010000000;
        samples[9] = 16'b1111111001110001;
        samples[10] = 16'b1111110100110011;
        samples[11] = 16'b1111110111011011;
        samples[12] = 16'b0000000110010010;
        samples[13] = 16'b0000010001100111;
        samples[14] = 16'b1111110011100001;
        samples[15] = 16'b1111111001111011;
        samples[16] = 16'b1111110111110001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000001100010;
        samples[1] = 16'b1111111101000110;
        samples[2] = 16'b1111111110100111;
        samples[3] = 16'b0000000000001011;
        samples[4] = 16'b0000000110010010;
        samples[5] = 16'b1111111101001001;
        samples[6] = 16'b1111111100000100;
        samples[7] = 16'b1111111101111011;
        samples[8] = 16'b0000010100010000;
        samples[9] = 16'b1111111010000111;
        samples[10] = 16'b1111110101001111;
        samples[11] = 16'b1111110100110110;
        samples[12] = 16'b0000001000000010;
        samples[13] = 16'b0000001011000001;
        samples[14] = 16'b1111101010110010;
        samples[15] = 16'b1111111010011010;
        samples[16] = 16'b1111111000110000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000001011100;
        samples[1] = 16'b1111111100100111;
        samples[2] = 16'b1111111111000011;
        samples[3] = 16'b1111111111001001;
        samples[4] = 16'b0000000100010101;
        samples[5] = 16'b1111111101011100;
        samples[6] = 16'b1111111101101100;
        samples[7] = 16'b1111111100110011;
        samples[8] = 16'b0000001111101101;
        samples[9] = 16'b1111110110101101;
        samples[10] = 16'b1111111010011101;
        samples[11] = 16'b1111110111010010;
        samples[12] = 16'b0000001001111100;
        samples[13] = 16'b1111110111011111;
        samples[14] = 16'b1111101101101010;
        samples[15] = 16'b1111111010100000;
        samples[16] = 16'b1111111010001010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000000010001;
        samples[1] = 16'b1111111100001110;
        samples[2] = 16'b1111111111101001;
        samples[3] = 16'b0000000000111010;
        samples[4] = 16'b0000000010010100;
        samples[5] = 16'b1111111101101000;
        samples[6] = 16'b1111111111000110;
        samples[7] = 16'b1111111110000101;
        samples[8] = 16'b0000001111000111;
        samples[9] = 16'b1111111100011101;
        samples[10] = 16'b1111111000110011;
        samples[11] = 16'b1111111000010111;
        samples[12] = 16'b0000001110010101;
        samples[13] = 16'b1111110111010010;
        samples[14] = 16'b1111101111100111;
        samples[15] = 16'b1111111011101000;
        samples[16] = 16'b1111111011100010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000000000010;
        samples[1] = 16'b1111111100010111;
        samples[2] = 16'b1111111111000110;
        samples[3] = 16'b0000000001101001;
        samples[4] = 16'b1111111111111110;
        samples[5] = 16'b1111111101000011;
        samples[6] = 16'b1111111111110010;
        samples[7] = 16'b0000000000011110;
        samples[8] = 16'b0000001010001111;
        samples[9] = 16'b1111111110101010;
        samples[10] = 16'b1111111001111110;
        samples[11] = 16'b1111111001111110;
        samples[12] = 16'b0000010001001000;
        samples[13] = 16'b0000000000010111;
        samples[14] = 16'b1111110011010101;
        samples[15] = 16'b1111111100011101;
        samples[16] = 16'b1111111100101010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111111100010;
        samples[1] = 16'b1111111100110110;
        samples[2] = 16'b1111111111001100;
        samples[3] = 16'b0000000000110100;
        samples[4] = 16'b1111111101101111;
        samples[5] = 16'b1111111100001011;
        samples[6] = 16'b0000000000111101;
        samples[7] = 16'b0000000001011111;
        samples[8] = 16'b0000000001010000;
        samples[9] = 16'b1111111110110011;
        samples[10] = 16'b1111111101001001;
        samples[11] = 16'b1111111100110110;
        samples[12] = 16'b0000011011101110;
        samples[13] = 16'b1111111111001001;
        samples[14] = 16'b1111111000100000;
        samples[15] = 16'b1111111100110011;
        samples[16] = 16'b1111111101111110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111111010110;
        samples[1] = 16'b1111111100010001;
        samples[2] = 16'b1111111111111011;
        samples[3] = 16'b0000000010111010;
        samples[4] = 16'b1111111100000001;
        samples[5] = 16'b1111111011011100;
        samples[6] = 16'b0000000011101001;
        samples[7] = 16'b0000000011011111;
        samples[8] = 16'b1111111000101010;
        samples[9] = 16'b0000000100001011;
        samples[10] = 16'b0000000011011001;
        samples[11] = 16'b0000000001101001;
        samples[12] = 16'b0000100000000100;
        samples[13] = 16'b0000010101000101;
        samples[14] = 16'b1111111000000111;
        samples[15] = 16'b1111111110110011;
        samples[16] = 16'b0000000000111101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111111011100;
        samples[1] = 16'b1111111100100001;
        samples[2] = 16'b1111111111111011;
        samples[3] = 16'b0000000100011011;
        samples[4] = 16'b1111111011101000;
        samples[5] = 16'b1111111010110011;
        samples[6] = 16'b0000000100011011;
        samples[7] = 16'b0000000101011101;
        samples[8] = 16'b1111110111010101;
        samples[9] = 16'b1111111111011111;
        samples[10] = 16'b0000000110101110;
        samples[11] = 16'b0000000100000010;
        samples[12] = 16'b0000100111101111;
        samples[13] = 16'b0000000100000101;
        samples[14] = 16'b1111111010001110;
        samples[15] = 16'b1111111111000110;
        samples[16] = 16'b0000000010011000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111111010011;
        samples[1] = 16'b1111111101101100;
        samples[2] = 16'b0000000001100010;
        samples[3] = 16'b0000000011100011;
        samples[4] = 16'b1111111100101010;
        samples[5] = 16'b1111111011100010;
        samples[6] = 16'b0000000100110111;
        samples[7] = 16'b0000000101000000;
        samples[8] = 16'b1111111101110010;
        samples[9] = 16'b1111111011111000;
        samples[10] = 16'b0000000101100110;
        samples[11] = 16'b0000000001011100;
        samples[12] = 16'b0000010010001001;
        samples[13] = 16'b0000000110101000;
        samples[14] = 16'b1111110011110111;
        samples[15] = 16'b1111111110110111;
        samples[16] = 16'b0000000001110010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000000101010;
        samples[1] = 16'b1111111110010001;
        samples[2] = 16'b0000000001101111;
        samples[3] = 16'b0000000100111101;
        samples[4] = 16'b1111111110101101;
        samples[5] = 16'b1111111101000011;
        samples[6] = 16'b0000000100001000;
        samples[7] = 16'b0000000101110010;
        samples[8] = 16'b0000000001001101;
        samples[9] = 16'b1111111110001110;
        samples[10] = 16'b0000000101110110;
        samples[11] = 16'b0000000010000010;
        samples[12] = 16'b0000000100101110;
        samples[13] = 16'b0000010001001000;
        samples[14] = 16'b1111110100110110;
        samples[15] = 16'b0000000000000101;
        samples[16] = 16'b0000000010101101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000010100111;
        samples[1] = 16'b1111111110011110;
        samples[2] = 16'b0000000000111101;
        samples[3] = 16'b0000000101110110;
        samples[4] = 16'b0000000000110111;
        samples[5] = 16'b1111111101011001;
        samples[6] = 16'b0000000011101100;
        samples[7] = 16'b0000000101111100;
        samples[8] = 16'b0000000000100001;
        samples[9] = 16'b0000000101101001;
        samples[10] = 16'b0000000010111010;
        samples[11] = 16'b0000000001101100;
        samples[12] = 16'b0000000110000010;
        samples[13] = 16'b0000000001010110;
        samples[14] = 16'b1111111000011010;
        samples[15] = 16'b0000000001011001;
        samples[16] = 16'b0000000011001101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101000000;
        samples[1] = 16'b1111111111000110;
        samples[2] = 16'b0000000001000000;
        samples[3] = 16'b0000000011101100;
        samples[4] = 16'b0000000011011001;
        samples[5] = 16'b1111111110001011;
        samples[6] = 16'b0000000011101001;
        samples[7] = 16'b0000000011110010;
        samples[8] = 16'b0000000011100110;
        samples[9] = 16'b0000001000100101;
        samples[10] = 16'b0000000000111101;
        samples[11] = 16'b1111111111111000;
        samples[12] = 16'b0000000101010011;
        samples[13] = 16'b0000010001100111;
        samples[14] = 16'b1111111000110000;
        samples[15] = 16'b0000000010011011;
        samples[16] = 16'b0000000011010110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101111001;
        samples[1] = 16'b1111111110101101;
        samples[2] = 16'b1111111111110101;
        samples[3] = 16'b0000000100110100;
        samples[4] = 16'b0000000100001011;
        samples[5] = 16'b1111111101001100;
        samples[6] = 16'b0000000010100100;
        samples[7] = 16'b0000000101010110;
        samples[8] = 16'b1111111010110011;
        samples[9] = 16'b0000001001011010;
        samples[10] = 16'b0000000110010101;
        samples[11] = 16'b0000000011110101;
        samples[12] = 16'b0000010100101111;
        samples[13] = 16'b0000001010010101;
        samples[14] = 16'b1111111100010100;
        samples[15] = 16'b0000000010101010;
        samples[16] = 16'b0000000011111100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110111010;
        samples[1] = 16'b1111111110110111;
        samples[2] = 16'b1111111110110011;
        samples[3] = 16'b0000000100100001;
        samples[4] = 16'b0000000101001101;
        samples[5] = 16'b1111111100101010;
        samples[6] = 16'b0000000001111111;
        samples[7] = 16'b0000000101010110;
        samples[8] = 16'b1111111000000111;
        samples[9] = 16'b0000001001000100;
        samples[10] = 16'b0000001001000001;
        samples[11] = 16'b0000000011101100;
        samples[12] = 16'b0000011010011101;
        samples[13] = 16'b1111111111111110;
        samples[14] = 16'b1111111011010101;
        samples[15] = 16'b0000000010101101;
        samples[16] = 16'b0000000100011110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000111011101;
        samples[1] = 16'b1111111111001100;
        samples[2] = 16'b1111111101010011;
        samples[3] = 16'b0000000011111000;
        samples[4] = 16'b0000000110011011;
        samples[5] = 16'b1111111011101110;
        samples[6] = 16'b0000000000110000;
        samples[7] = 16'b0000000100111010;
        samples[8] = 16'b0000000011010011;
        samples[9] = 16'b0000000000100001;
        samples[10] = 16'b0000000100101011;
        samples[11] = 16'b0000000010000101;
        samples[12] = 16'b0000000111111001;
        samples[13] = 16'b0000001000101000;
        samples[14] = 16'b1111111101110101;
        samples[15] = 16'b0000000000110000;
        samples[16] = 16'b0000000010011110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000111111111;
        samples[1] = 16'b0000000000010001;
        samples[2] = 16'b1111111101001100;
        samples[3] = 16'b0000000011101001;
        samples[4] = 16'b0000000111110011;
        samples[5] = 16'b1111111100100111;
        samples[6] = 16'b0000000000000010;
        samples[7] = 16'b0000000100100100;
        samples[8] = 16'b0000000110101110;
        samples[9] = 16'b0000000010011110;
        samples[10] = 16'b0000000011010110;
        samples[11] = 16'b0000000001100010;
        samples[12] = 16'b0000000001101111;
        samples[13] = 16'b0000000101111100;
        samples[14] = 16'b1111111100100100;
        samples[15] = 16'b0000000001001001;
        samples[16] = 16'b0000000001111011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000001000011110;
        samples[1] = 16'b0000000000110100;
        samples[2] = 16'b1111111100100111;
        samples[3] = 16'b0000000011100110;
        samples[4] = 16'b0000000111111111;
        samples[5] = 16'b1111111101011111;
        samples[6] = 16'b1111111111111011;
        samples[7] = 16'b0000000100001000;
        samples[8] = 16'b0000000101010011;
        samples[9] = 16'b0000000101000111;
        samples[10] = 16'b0000000100101110;
        samples[11] = 16'b0000000010100001;
        samples[12] = 16'b0000000000110000;
        samples[13] = 16'b0000000010011000;
        samples[14] = 16'b1111111101001100;
        samples[15] = 16'b0000000001110101;
        samples[16] = 16'b0000000010010100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000001000001100;
        samples[1] = 16'b0000000001100110;
        samples[2] = 16'b1111111100011101;
        samples[3] = 16'b0000000010001011;
        samples[4] = 16'b0000000111011101;
        samples[5] = 16'b1111111110000001;
        samples[6] = 16'b0000000000000101;
        samples[7] = 16'b0000000010110111;
        samples[8] = 16'b0000000110110111;
        samples[9] = 16'b0000000110000101;
        samples[10] = 16'b0000000001100110;
        samples[11] = 16'b0000000000010100;
        samples[12] = 16'b1111111100110000;
        samples[13] = 16'b0000011010001101;
        samples[14] = 16'b1111111111000011;
        samples[15] = 16'b0000000001011100;
        samples[16] = 16'b0000000001100110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000111001010;
        samples[1] = 16'b0000000010011110;
        samples[2] = 16'b1111111101000110;
        samples[3] = 16'b0000000001101001;
        samples[4] = 16'b0000000110001111;
        samples[5] = 16'b1111111110111101;
        samples[6] = 16'b0000000000001011;
        samples[7] = 16'b0000000011000000;
        samples[8] = 16'b0000000000011011;
        samples[9] = 16'b0000000011011001;
        samples[10] = 16'b0000000111011010;
        samples[11] = 16'b0000000001001001;
        samples[12] = 16'b0000010111100100;
        samples[13] = 16'b0000001111110110;
        samples[14] = 16'b1111111111111011;
        samples[15] = 16'b0000000000111010;
        samples[16] = 16'b0000000010101010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101010000;
        samples[1] = 16'b0000000001101001;
        samples[2] = 16'b1111111100010111;
        samples[3] = 16'b0000000011100110;
        samples[4] = 16'b0000000011110101;
        samples[5] = 16'b1111111110100001;
        samples[6] = 16'b0000000000000010;
        samples[7] = 16'b0000000100101110;
        samples[8] = 16'b1111110111010101;
        samples[9] = 16'b1111111111010000;
        samples[10] = 16'b0000001011111111;
        samples[11] = 16'b0000000110001011;
        samples[12] = 16'b0000011100110011;
        samples[13] = 16'b0000010000110010;
        samples[14] = 16'b0000000110100001;
        samples[15] = 16'b1111111111110010;
        samples[16] = 16'b0000000011110010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011010011;
        samples[1] = 16'b0000000000110100;
        samples[2] = 16'b1111111011111110;
        samples[3] = 16'b0000000100111101;
        samples[4] = 16'b0000000010000101;
        samples[5] = 16'b1111111101111011;
        samples[6] = 16'b1111111111110010;
        samples[7] = 16'b0000000101010110;
        samples[8] = 16'b1111111100110011;
        samples[9] = 16'b1111111001010101;
        samples[10] = 16'b0000001000100001;
        samples[11] = 16'b0000000110000101;
        samples[12] = 16'b0000011101000101;
        samples[13] = 16'b0000000101101001;
        samples[14] = 16'b0000000111101111;
        samples[15] = 16'b1111111110001011;
        samples[16] = 16'b0000000011001101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000000111010;
        samples[1] = 16'b0000000001010011;
        samples[2] = 16'b1111111100011101;
        samples[3] = 16'b0000000101011001;
        samples[4] = 16'b1111111111110010;
        samples[5] = 16'b1111111110010111;
        samples[6] = 16'b1111111111010000;
        samples[7] = 16'b0000000110110100;
        samples[8] = 16'b1111111010110110;
        samples[9] = 16'b1111111110100100;
        samples[10] = 16'b0000000111101100;
        samples[11] = 16'b0000000010101010;
        samples[12] = 16'b0000011001100001;
        samples[13] = 16'b1111111011011111;
        samples[14] = 16'b0000000001101001;
        samples[15] = 16'b1111111110110111;
        samples[16] = 16'b0000000010011011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111111001100;
        samples[1] = 16'b0000000001101100;
        samples[2] = 16'b1111111100000100;
        samples[3] = 16'b0000000110101011;
        samples[4] = 16'b1111111110100111;
        samples[5] = 16'b1111111110011010;
        samples[6] = 16'b1111111110110000;
        samples[7] = 16'b0000000111111001;
        samples[8] = 16'b1111111101001100;
        samples[9] = 16'b0000000010000010;
        samples[10] = 16'b0000000100011000;
        samples[11] = 16'b1111111111111011;
        samples[12] = 16'b0000010100111011;
        samples[13] = 16'b1111101110011111;
        samples[14] = 16'b1111111010000111;
        samples[15] = 16'b1111111111101001;
        samples[16] = 16'b0000000001011111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110101101;
        samples[1] = 16'b0000000001101001;
        samples[2] = 16'b1111111100011101;
        samples[3] = 16'b0000000011101100;
        samples[4] = 16'b1111111110001110;
        samples[5] = 16'b1111111111010000;
        samples[6] = 16'b1111111111101001;
        samples[7] = 16'b0000000011011100;
        samples[8] = 16'b0000000001011100;
        samples[9] = 16'b0000000011111100;
        samples[10] = 16'b0000000000011011;
        samples[11] = 16'b1111111100001000;
        samples[12] = 16'b0000001010000101;
        samples[13] = 16'b1111110111101110;
        samples[14] = 16'b1111111001111110;
        samples[15] = 16'b0000000000010111;
        samples[16] = 16'b0000000000110100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101111000;
        samples[1] = 16'b0000000001100110;
        samples[2] = 16'b1111111011101000;
        samples[3] = 16'b0000000011101111;
        samples[4] = 16'b1111111101010110;
        samples[5] = 16'b1111111111111011;
        samples[6] = 16'b1111111111000000;
        samples[7] = 16'b0000000010100111;
        samples[8] = 16'b0000000101000100;
        samples[9] = 16'b0000000001111000;
        samples[10] = 16'b1111111101110101;
        samples[11] = 16'b1111111010010100;
        samples[12] = 16'b0000000110000101;
        samples[13] = 16'b1111111011001100;
        samples[14] = 16'b1111111010101010;
        samples[15] = 16'b1111111111110010;
        samples[16] = 16'b1111111111110101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111111010110;
        samples[1] = 16'b0000000010101010;
        samples[2] = 16'b1111111011101110;
        samples[3] = 16'b0000000000011011;
        samples[4] = 16'b1111111110100111;
        samples[5] = 16'b0000000001110101;
        samples[6] = 16'b1111111101101111;
        samples[7] = 16'b0000000000000010;
        samples[8] = 16'b0000000010010001;
        samples[9] = 16'b1111111111011001;
        samples[10] = 16'b0000000000111010;
        samples[11] = 16'b1111111011001001;
        samples[12] = 16'b0000010110001010;
        samples[13] = 16'b1111110010010000;
        samples[14] = 16'b1111111101111110;
        samples[15] = 16'b1111111111010110;
        samples[16] = 16'b0000000000000010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110110000;
        samples[1] = 16'b0000000001000110;
        samples[2] = 16'b1111111001011100;
        samples[3] = 16'b0000000001111011;
        samples[4] = 16'b1111111100110011;
        samples[5] = 16'b0000000001001001;
        samples[6] = 16'b1111111011101110;
        samples[7] = 16'b0000000001100010;
        samples[8] = 16'b1111111100001110;
        samples[9] = 16'b1111111110100111;
        samples[10] = 16'b0000000001100010;
        samples[11] = 16'b1111111110111101;
        samples[12] = 16'b0000000110101011;
        samples[13] = 16'b1111111000010001;
        samples[14] = 16'b0000000101000111;
        samples[15] = 16'b1111111110100111;
        samples[16] = 16'b0000000000000010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110100111;
        samples[1] = 16'b0000000000100100;
        samples[2] = 16'b1111111001011111;
        samples[3] = 16'b0000000010111101;
        samples[4] = 16'b1111111100110000;
        samples[5] = 16'b0000000001011001;
        samples[6] = 16'b1111111011000110;
        samples[7] = 16'b0000000010010100;
        samples[8] = 16'b1111111111000011;
        samples[9] = 16'b1111111110011110;
        samples[10] = 16'b1111111111011111;
        samples[11] = 16'b1111111101100010;
        samples[12] = 16'b1111111001001111;
        samples[13] = 16'b1111111100001011;
        samples[14] = 16'b0000000010001011;
        samples[15] = 16'b1111111110000101;
        samples[16] = 16'b1111111111101111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110111010;
        samples[1] = 16'b0000000000100100;
        samples[2] = 16'b1111111001100101;
        samples[3] = 16'b0000000001011100;
        samples[4] = 16'b1111111101101111;
        samples[5] = 16'b0000000001001001;
        samples[6] = 16'b1111111010100111;
        samples[7] = 16'b0000000001000000;
        samples[8] = 16'b1111111101100101;
        samples[9] = 16'b1111111100011101;
        samples[10] = 16'b0000000000001110;
        samples[11] = 16'b1111111101110010;
        samples[12] = 16'b0000000111000111;
        samples[13] = 16'b1111110100100110;
        samples[14] = 16'b0000000010000010;
        samples[15] = 16'b1111111101001100;
        samples[16] = 16'b1111111110101101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111111000000;
        samples[1] = 16'b0000000000011110;
        samples[2] = 16'b1111111001101000;
        samples[3] = 16'b0000000000001011;
        samples[4] = 16'b1111111110100100;
        samples[5] = 16'b0000000000111101;
        samples[6] = 16'b1111111010010001;
        samples[7] = 16'b1111111111011100;
        samples[8] = 16'b1111111111011001;
        samples[9] = 16'b1111111011011100;
        samples[10] = 16'b1111111111000000;
        samples[11] = 16'b1111111110110111;
        samples[12] = 16'b1111111001101000;
        samples[13] = 16'b0000010000110010;
        samples[14] = 16'b0000000011100011;
        samples[15] = 16'b1111111101001001;
        samples[16] = 16'b1111111101100101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101101000;
        samples[1] = 16'b1111111111000011;
        samples[2] = 16'b1111111001011000;
        samples[3] = 16'b0000000000110100;
        samples[4] = 16'b1111111110100001;
        samples[5] = 16'b0000000000001000;
        samples[6] = 16'b1111111001100010;
        samples[7] = 16'b1111111110101010;
        samples[8] = 16'b0000001000110100;
        samples[9] = 16'b1111110011001111;
        samples[10] = 16'b1111111000110000;
        samples[11] = 16'b1111111011101011;
        samples[12] = 16'b0000000001111111;
        samples[13] = 16'b0000000101111001;
        samples[14] = 16'b0000000010110001;
        samples[15] = 16'b1111111010101101;
        samples[16] = 16'b1111111011100010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101101000;
        samples[1] = 16'b1111111111101100;
        samples[2] = 16'b1111111010001010;
        samples[3] = 16'b1111111101110010;
        samples[4] = 16'b1111111110110000;
        samples[5] = 16'b0000000000100001;
        samples[6] = 16'b1111111001111110;
        samples[7] = 16'b1111111011111011;
        samples[8] = 16'b0000000011000000;
        samples[9] = 16'b1111110000001101;
        samples[10] = 16'b1111111110001110;
        samples[11] = 16'b1111111010100111;
        samples[12] = 16'b0000010000000000;
        samples[13] = 16'b1111111111101111;
        samples[14] = 16'b0000000001001001;
        samples[15] = 16'b1111111010001010;
        samples[16] = 16'b1111111011100101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101000110;
        samples[1] = 16'b1111111111000011;
        samples[2] = 16'b1111111010000001;
        samples[3] = 16'b1111111110110000;
        samples[4] = 16'b1111111110101010;
        samples[5] = 16'b0000000000000101;
        samples[6] = 16'b1111111001101000;
        samples[7] = 16'b1111111100011010;
        samples[8] = 16'b0000000111000100;
        samples[9] = 16'b1111101111100001;
        samples[10] = 16'b1111111100000100;
        samples[11] = 16'b1111111100111010;
        samples[12] = 16'b0000001011010111;
        samples[13] = 16'b0000000001101001;
        samples[14] = 16'b0000000101010000;
        samples[15] = 16'b1111111010010001;
        samples[16] = 16'b1111111011001001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011100101;
        samples[1] = 16'b1111111101101100;
        samples[2] = 16'b1111111001010010;
        samples[3] = 16'b0000000001101001;
        samples[4] = 16'b1111111101101111;
        samples[5] = 16'b1111111111010110;
        samples[6] = 16'b1111111001001111;
        samples[7] = 16'b1111111101111000;
        samples[8] = 16'b0000000010101010;
        samples[9] = 16'b1111110110100110;
        samples[10] = 16'b1111111001111000;
        samples[11] = 16'b1111111100100100;
        samples[12] = 16'b0000000000100111;
        samples[13] = 16'b1111011110001111;
        samples[14] = 16'b0000000100111101;
        samples[15] = 16'b1111111010100111;
        samples[16] = 16'b1111111011001100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011101110;
        samples[1] = 16'b1111111111010011;
        samples[2] = 16'b1111111010110000;
        samples[3] = 16'b1111111111001001;
        samples[4] = 16'b1111111110011110;
        samples[5] = 16'b0000000000010111;
        samples[6] = 16'b1111111010010001;
        samples[7] = 16'b1111111011101110;
        samples[8] = 16'b1111111101001111;
        samples[9] = 16'b1111111101110010;
        samples[10] = 16'b1111111100101010;
        samples[11] = 16'b1111111000100110;
        samples[12] = 16'b0000000011110010;
        samples[13] = 16'b1111011110000010;
        samples[14] = 16'b1111111100101101;
        samples[15] = 16'b1111111011001100;
        samples[16] = 16'b1111111011111110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111010110011;
        samples[1] = 16'b1111111111110101;
        samples[2] = 16'b1111111011011111;
        samples[3] = 16'b1111111110111101;
        samples[4] = 16'b1111111110110011;
        samples[5] = 16'b0000000000001000;
        samples[6] = 16'b1111111010001010;
        samples[7] = 16'b1111111011111011;
        samples[8] = 16'b0000000011100011;
        samples[9] = 16'b1111111100010100;
        samples[10] = 16'b1111111000100000;
        samples[11] = 16'b1111111000000100;
        samples[12] = 16'b1111110111011000;
        samples[13] = 16'b1111111010010001;
        samples[14] = 16'b1111111011100101;
        samples[15] = 16'b1111111001111000;
        samples[16] = 16'b1111111011000000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111010101101;
        samples[1] = 16'b1111111111111011;
        samples[2] = 16'b1111111100001000;
        samples[3] = 16'b1111111110110111;
        samples[4] = 16'b1111111111010011;
        samples[5] = 16'b1111111111011100;
        samples[6] = 16'b1111111011001100;
        samples[7] = 16'b1111111011101110;
        samples[8] = 16'b1111111111110010;
        samples[9] = 16'b1111111101100010;
        samples[10] = 16'b1111111000001010;
        samples[11] = 16'b1111111010000100;
        samples[12] = 16'b0000000010111101;
        samples[13] = 16'b1111110010100110;
        samples[14] = 16'b1111111101110010;
        samples[15] = 16'b1111111001000011;
        samples[16] = 16'b1111111011010101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111010100111;
        samples[1] = 16'b1111111111101001;
        samples[2] = 16'b1111111101101111;
        samples[3] = 16'b1111111101010110;
        samples[4] = 16'b1111111110111010;
        samples[5] = 16'b1111111110101101;
        samples[6] = 16'b1111111100110011;
        samples[7] = 16'b1111111010111001;
        samples[8] = 16'b1111111110110000;
        samples[9] = 16'b1111110111111000;
        samples[10] = 16'b1111111011110010;
        samples[11] = 16'b1111111011000011;
        samples[12] = 16'b0000000111000001;
        samples[13] = 16'b1111111101000011;
        samples[14] = 16'b1111111011000000;
        samples[15] = 16'b1111110111101000;
        samples[16] = 16'b1111111011110101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111000111001;
        samples[1] = 16'b0000000000001011;
        samples[2] = 16'b1111111111010011;
        samples[3] = 16'b1111111101000000;
        samples[4] = 16'b1111111101101111;
        samples[5] = 16'b1111111101000110;
        samples[6] = 16'b1111111101000011;
        samples[7] = 16'b1111111101011111;
        samples[8] = 16'b0000000100001110;
        samples[9] = 16'b1111101100100010;
        samples[10] = 16'b1111111011000000;
        samples[11] = 16'b1111111100010100;
        samples[12] = 16'b0000000110101110;
        samples[13] = 16'b1111111110001110;
        samples[14] = 16'b1111111001000011;
        samples[15] = 16'b1111110100111100;
        samples[16] = 16'b1111111010011010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111001100;
        samples[1] = 16'b1111111111111110;
        samples[2] = 16'b1111111111101001;
        samples[3] = 16'b1111111111000110;
        samples[4] = 16'b1111111100100001;
        samples[5] = 16'b1111111011110010;
        samples[6] = 16'b1111111101100101;
        samples[7] = 16'b1111111111111110;
        samples[8] = 16'b0000000100111010;
        samples[9] = 16'b1111101101111101;
        samples[10] = 16'b1111111000010001;
        samples[11] = 16'b1111111100101101;
        samples[12] = 16'b1111111111101100;
        samples[13] = 16'b1111110110110110;
        samples[14] = 16'b1111111011011111;
        samples[15] = 16'b1111110100100110;
        samples[16] = 16'b1111111010010100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111001001;
        samples[1] = 16'b1111111111110010;
        samples[2] = 16'b0000000000100001;
        samples[3] = 16'b1111111110010001;
        samples[4] = 16'b1111111100011010;
        samples[5] = 16'b1111111100100111;
        samples[6] = 16'b1111111111000000;
        samples[7] = 16'b1111111101101000;
        samples[8] = 16'b0000000011011001;
        samples[9] = 16'b1111110011001111;
        samples[10] = 16'b1111111000100000;
        samples[11] = 16'b1111111000011010;
        samples[12] = 16'b0000000111010000;
        samples[13] = 16'b1111101010011100;
        samples[14] = 16'b1111110100011010;
        samples[15] = 16'b1111110101000101;
        samples[16] = 16'b1111111011011111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111000110;
        samples[1] = 16'b1111111111101111;
        samples[2] = 16'b0000000000110000;
        samples[3] = 16'b1111111110110011;
        samples[4] = 16'b1111111100010001;
        samples[5] = 16'b1111111101011001;
        samples[6] = 16'b1111111111001001;
        samples[7] = 16'b1111111101100101;
        samples[8] = 16'b0000001100010101;
        samples[9] = 16'b1111110010110010;
        samples[10] = 16'b1111110010000111;
        samples[11] = 16'b1111110110110011;
        samples[12] = 16'b0000000110001000;
        samples[13] = 16'b1111110100010000;
        samples[14] = 16'b1111110110000001;
        samples[15] = 16'b1111110011100001;
        samples[16] = 16'b1111111011001100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111100101;
        samples[1] = 16'b1111111111111011;
        samples[2] = 16'b0000000000000010;
        samples[3] = 16'b1111111110101010;
        samples[4] = 16'b1111111011101011;
        samples[5] = 16'b1111111101111110;
        samples[6] = 16'b1111111110100100;
        samples[7] = 16'b1111111110000001;
        samples[8] = 16'b0000001000101000;
        samples[9] = 16'b1111110101100101;
        samples[10] = 16'b1111110001011011;
        samples[11] = 16'b1111111000100011;
        samples[12] = 16'b0000000100110111;
        samples[13] = 16'b0000000010000101;
        samples[14] = 16'b1111111000111111;
        samples[15] = 16'b1111110011101110;
        samples[16] = 16'b1111111011101011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111101110;
        samples[1] = 16'b1111111111000011;
        samples[2] = 16'b1111111111011111;
        samples[3] = 16'b1111111110101010;
        samples[4] = 16'b1111111010000111;
        samples[5] = 16'b1111111101111110;
        samples[6] = 16'b1111111110010111;
        samples[7] = 16'b1111111110100001;
        samples[8] = 16'b0000000010001000;
        samples[9] = 16'b1111110001011000;
        samples[10] = 16'b1111110110000100;
        samples[11] = 16'b1111111001111110;
        samples[12] = 16'b0000011100110000;
        samples[13] = 16'b1111101000000011;
        samples[14] = 16'b1111110110111100;
        samples[15] = 16'b1111110011000010;
        samples[16] = 16'b1111111100010111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111000001101;
        samples[1] = 16'b1111111110101101;
        samples[2] = 16'b1111111111101100;
        samples[3] = 16'b1111111110000001;
        samples[4] = 16'b1111111000101010;
        samples[5] = 16'b1111111110010001;
        samples[6] = 16'b1111111111000011;
        samples[7] = 16'b1111111110101101;
        samples[8] = 16'b1111111111001100;
        samples[9] = 16'b1111101111101010;
        samples[10] = 16'b1111111001100010;
        samples[11] = 16'b1111111010010001;
        samples[12] = 16'b0000010100100010;
        samples[13] = 16'b0000000000101101;
        samples[14] = 16'b1111110101000010;
        samples[15] = 16'b1111110011011000;
        samples[16] = 16'b1111111100110000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111111011;
        samples[1] = 16'b1111111110000101;
        samples[2] = 16'b1111111111000011;
        samples[3] = 16'b1111111111000000;
        samples[4] = 16'b1111110111101000;
        samples[5] = 16'b1111111101111110;
        samples[6] = 16'b1111111110001110;
        samples[7] = 16'b0000000000000101;
        samples[8] = 16'b0000000011000000;
        samples[9] = 16'b1111101000001001;
        samples[10] = 16'b1111111010000111;
        samples[11] = 16'b1111111011100101;
        samples[12] = 16'b0000000110110100;
        samples[13] = 16'b0000000000000101;
        samples[14] = 16'b1111110101001001;
        samples[15] = 16'b1111110010110010;
        samples[16] = 16'b1111111011011111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111110100;
        samples[1] = 16'b1111111101001001;
        samples[2] = 16'b1111111110110000;
        samples[3] = 16'b0000000000100100;
        samples[4] = 16'b1111110111011000;
        samples[5] = 16'b1111111110011010;
        samples[6] = 16'b1111111101111011;
        samples[7] = 16'b0000000000100111;
        samples[8] = 16'b0000000111100011;
        samples[9] = 16'b1111101011110111;
        samples[10] = 16'b1111110110100110;
        samples[11] = 16'b1111111001011100;
        samples[12] = 16'b1111110100111001;
        samples[13] = 16'b1111110100111100;
        samples[14] = 16'b1111110100000100;
        samples[15] = 16'b1111110011100100;
        samples[16] = 16'b1111111010111100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111000101010;
        samples[1] = 16'b1111111101101000;
        samples[2] = 16'b1111111110111101;
        samples[3] = 16'b1111111111011100;
        samples[4] = 16'b1111111000011101;
        samples[5] = 16'b1111111111000110;
        samples[6] = 16'b1111111110100111;
        samples[7] = 16'b1111111110100111;
        samples[8] = 16'b0000001101000111;
        samples[9] = 16'b1111101101100001;
        samples[10] = 16'b1111110011000010;
        samples[11] = 16'b1111110101110111;
        samples[12] = 16'b1111111100010001;
        samples[13] = 16'b1111110011100100;
        samples[14] = 16'b1111110001111101;
        samples[15] = 16'b1111110011001111;
        samples[16] = 16'b1111111010011010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111000011101;
        samples[1] = 16'b1111111101101100;
        samples[2] = 16'b1111111110000001;
        samples[3] = 16'b0000000001000000;
        samples[4] = 16'b1111110111110001;
        samples[5] = 16'b1111111110011010;
        samples[6] = 16'b1111111110001110;
        samples[7] = 16'b0000000000101010;
        samples[8] = 16'b0000001010001001;
        samples[9] = 16'b1111101011101101;
        samples[10] = 16'b1111110110000100;
        samples[11] = 16'b1111110111111000;
        samples[12] = 16'b1111111110111010;
        samples[13] = 16'b1111101100010011;
        samples[14] = 16'b1111110100110000;
        samples[15] = 16'b1111110010100000;
        samples[16] = 16'b1111111010111100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111000000100;
        samples[1] = 16'b1111111101011001;
        samples[2] = 16'b1111111101011001;
        samples[3] = 16'b0000000010110100;
        samples[4] = 16'b1111110111110001;
        samples[5] = 16'b1111111101110010;
        samples[6] = 16'b1111111110001000;
        samples[7] = 16'b0000000010001000;
        samples[8] = 16'b0000000111110011;
        samples[9] = 16'b1111101110000011;
        samples[10] = 16'b1111110100000001;
        samples[11] = 16'b1111111010111100;
        samples[12] = 16'b0000000001000110;
        samples[13] = 16'b1111101010110010;
        samples[14] = 16'b1111111001110001;
        samples[15] = 16'b1111110001110111;
        samples[16] = 16'b1111111011100101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111000101101;
        samples[1] = 16'b1111111101000000;
        samples[2] = 16'b1111111110010100;
        samples[3] = 16'b0000000001000000;
        samples[4] = 16'b1111110111111011;
        samples[5] = 16'b1111111110001000;
        samples[6] = 16'b1111111111011111;
        samples[7] = 16'b1111111111100010;
        samples[8] = 16'b0000000000011011;
        samples[9] = 16'b1111110001011110;
        samples[10] = 16'b1111111001001001;
        samples[11] = 16'b1111111011110101;
        samples[12] = 16'b0000010111010001;
        samples[13] = 16'b1111101011010001;
        samples[14] = 16'b1111110111010101;
        samples[15] = 16'b1111110001110111;
        samples[16] = 16'b1111111101011111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111111000;
        samples[1] = 16'b1111111011011100;
        samples[2] = 16'b1111111101101100;
        samples[3] = 16'b0000000011111100;
        samples[4] = 16'b1111110110101001;
        samples[5] = 16'b1111111101010110;
        samples[6] = 16'b1111111110010111;
        samples[7] = 16'b0000000010100100;
        samples[8] = 16'b1111111011001001;
        samples[9] = 16'b1111110011111010;
        samples[10] = 16'b1111111011011001;
        samples[11] = 16'b1111111100110000;
        samples[12] = 16'b1111110110011010;
        samples[13] = 16'b0000001101010111;
        samples[14] = 16'b1111110011111010;
        samples[15] = 16'b1111110001101011;
        samples[16] = 16'b1111111110001011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111010101;
        samples[1] = 16'b1111111011110010;
        samples[2] = 16'b1111111101100101;
        samples[3] = 16'b0000000011011100;
        samples[4] = 16'b1111110110111111;
        samples[5] = 16'b1111111101000000;
        samples[6] = 16'b1111111110001000;
        samples[7] = 16'b0000000010000010;
        samples[8] = 16'b1111111101010110;
        samples[9] = 16'b1111110001100001;
        samples[10] = 16'b1111111011010101;
        samples[11] = 16'b1111111100110011;
        samples[12] = 16'b1111111101101100;
        samples[13] = 16'b0000010100001101;
        samples[14] = 16'b1111110010101111;
        samples[15] = 16'b1111110001010010;
        samples[16] = 16'b1111111110101010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111110111111000;
        samples[1] = 16'b1111111010100011;
        samples[2] = 16'b1111111101000110;
        samples[3] = 16'b0000000011011111;
        samples[4] = 16'b1111110111001111;
        samples[5] = 16'b1111111011111011;
        samples[6] = 16'b1111111111000000;
        samples[7] = 16'b0000000000111010;
        samples[8] = 16'b1111111101110101;
        samples[9] = 16'b1111110010010110;
        samples[10] = 16'b1111111001110001;
        samples[11] = 16'b1111111111000110;
        samples[12] = 16'b1111110101011011;
        samples[13] = 16'b0000000010111010;
        samples[14] = 16'b1111110110010111;
        samples[15] = 16'b1111110001101011;
        samples[16] = 16'b1111111111011100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111000001101;
        samples[1] = 16'b1111111010110000;
        samples[2] = 16'b1111111100110000;
        samples[3] = 16'b0000000101000111;
        samples[4] = 16'b1111110111100010;
        samples[5] = 16'b1111111011001001;
        samples[6] = 16'b1111111111110010;
        samples[7] = 16'b0000000010010100;
        samples[8] = 16'b1111111001100101;
        samples[9] = 16'b1111111000010100;
        samples[10] = 16'b1111111001111000;
        samples[11] = 16'b0000000001010011;
        samples[12] = 16'b0000000011001101;
        samples[13] = 16'b1111110100100110;
        samples[14] = 16'b1111110111101110;
        samples[15] = 16'b1111110011011110;
        samples[16] = 16'b0000000001000011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111000110000;
        samples[1] = 16'b1111111100111101;
        samples[2] = 16'b1111111101101111;
        samples[3] = 16'b0000000010110001;
        samples[4] = 16'b1111111000000001;
        samples[5] = 16'b1111111011011100;
        samples[6] = 16'b0000000000110111;
        samples[7] = 16'b0000000001101111;
        samples[8] = 16'b1111111100001000;
        samples[9] = 16'b1111110110110000;
        samples[10] = 16'b1111111010100011;
        samples[11] = 16'b0000000000111101;
        samples[12] = 16'b1111111101101111;
        samples[13] = 16'b0000000000001011;
        samples[14] = 16'b1111111001010010;
        samples[15] = 16'b1111110100110110;
        samples[16] = 16'b0000000001011100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111001010101;
        samples[1] = 16'b1111111110001000;
        samples[2] = 16'b1111111110101010;
        samples[3] = 16'b0000000001101111;
        samples[4] = 16'b1111110111110001;
        samples[5] = 16'b1111111100110110;
        samples[6] = 16'b0000000001101100;
        samples[7] = 16'b0000000001011111;
        samples[8] = 16'b1111111010110110;
        samples[9] = 16'b1111111000110011;
        samples[10] = 16'b1111111011000000;
        samples[11] = 16'b0000000001001101;
        samples[12] = 16'b0000001000000010;
        samples[13] = 16'b1111101011011010;
        samples[14] = 16'b1111111010000100;
        samples[15] = 16'b1111110110110000;
        samples[16] = 16'b0000000010011110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111010100011;
        samples[1] = 16'b1111111110110011;
        samples[2] = 16'b1111111110100001;
        samples[3] = 16'b0000000010101101;
        samples[4] = 16'b1111110111110001;
        samples[5] = 16'b1111111110111010;
        samples[6] = 16'b0000000010100001;
        samples[7] = 16'b0000000001010011;
        samples[8] = 16'b1111110111110001;
        samples[9] = 16'b1111111101011111;
        samples[10] = 16'b1111111110010100;
        samples[11] = 16'b0000000001101001;
        samples[12] = 16'b1111111110010001;
        samples[13] = 16'b0000010000101000;
        samples[14] = 16'b1111111100100100;
        samples[15] = 16'b1111111001111110;
        samples[16] = 16'b0000000100010010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111011100101;
        samples[1] = 16'b0000000000000010;
        samples[2] = 16'b1111111110110111;
        samples[3] = 16'b0000000001111111;
        samples[4] = 16'b1111111000000001;
        samples[5] = 16'b0000000001000000;
        samples[6] = 16'b0000000011000000;
        samples[7] = 16'b0000000000001110;
        samples[8] = 16'b1111111101100010;
        samples[9] = 16'b1111111011101110;
        samples[10] = 16'b1111111101101100;
        samples[11] = 16'b0000000000000010;
        samples[12] = 16'b1111111001011111;
        samples[13] = 16'b0000011110000111;
        samples[14] = 16'b1111111011100101;
        samples[15] = 16'b1111111100000001;
        samples[16] = 16'b0000000100100100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101001111;
        samples[1] = 16'b0000000000111101;
        samples[2] = 16'b1111111110001000;
        samples[3] = 16'b0000000001101100;
        samples[4] = 16'b1111111000110110;
        samples[5] = 16'b0000000010001000;
        samples[6] = 16'b0000000010011110;
        samples[7] = 16'b0000000000011011;
        samples[8] = 16'b1111111001001111;
        samples[9] = 16'b1111111011111000;
        samples[10] = 16'b0000000001000000;
        samples[11] = 16'b0000000011011100;
        samples[12] = 16'b0000001100011111;
        samples[13] = 16'b0000000000001000;
        samples[14] = 16'b0000000000001110;
        samples[15] = 16'b1111111110001110;
        samples[16] = 16'b0000000100110111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110111101;
        samples[1] = 16'b0000000000110111;
        samples[2] = 16'b1111111101101000;
        samples[3] = 16'b0000000001111000;
        samples[4] = 16'b1111111001011000;
        samples[5] = 16'b0000000010111010;
        samples[6] = 16'b0000000010100001;
        samples[7] = 16'b0000000000100100;
        samples[8] = 16'b1111110100100000;
        samples[9] = 16'b0000000011100110;
        samples[10] = 16'b0000000000110000;
        samples[11] = 16'b0000000011010000;
        samples[12] = 16'b0000000100000010;
        samples[13] = 16'b1111101110111000;
        samples[14] = 16'b0000000000000010;
        samples[15] = 16'b0000000001000011;
        samples[16] = 16'b0000000101011101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000000010001;
        samples[1] = 16'b0000000001111000;
        samples[2] = 16'b1111111110001110;
        samples[3] = 16'b0000000001100110;
        samples[4] = 16'b1111111010000001;
        samples[5] = 16'b0000000011101111;
        samples[6] = 16'b0000000011000011;
        samples[7] = 16'b0000000001000110;
        samples[8] = 16'b1111110100000100;
        samples[9] = 16'b0000001001011010;
        samples[10] = 16'b0000000001010000;
        samples[11] = 16'b0000000010011011;
        samples[12] = 16'b1111111111111000;
        samples[13] = 16'b1111110001010010;
        samples[14] = 16'b1111111011110010;
        samples[15] = 16'b0000000011110010;
        samples[16] = 16'b0000000110011110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000010001011;
        samples[1] = 16'b0000000001011100;
        samples[2] = 16'b1111111110101101;
        samples[3] = 16'b0000000000001110;
        samples[4] = 16'b1111111010011101;
        samples[5] = 16'b0000000011111000;
        samples[6] = 16'b0000000011011001;
        samples[7] = 16'b0000000000110100;
        samples[8] = 16'b1111101010110101;
        samples[9] = 16'b0000001011101101;
        samples[10] = 16'b0000001000000101;
        samples[11] = 16'b0000000101101001;
        samples[12] = 16'b0000000110100100;
        samples[13] = 16'b1111110100001101;
        samples[14] = 16'b1111111101001111;
        samples[15] = 16'b0000000101101111;
        samples[16] = 16'b0000000111000111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011010011;
        samples[1] = 16'b0000000000110111;
        samples[2] = 16'b1111111111111011;
        samples[3] = 16'b0000000000110000;
        samples[4] = 16'b1111111011000011;
        samples[5] = 16'b0000000100011011;
        samples[6] = 16'b0000000011110010;
        samples[7] = 16'b0000000001101001;
        samples[8] = 16'b1111101011101101;
        samples[9] = 16'b0000001101000111;
        samples[10] = 16'b0000000111100110;
        samples[11] = 16'b0000000111011010;
        samples[12] = 16'b0000000110001011;
        samples[13] = 16'b1111110010110010;
        samples[14] = 16'b1111111111001100;
        samples[15] = 16'b0000000111100011;
        samples[16] = 16'b0000000111011101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011010000;
        samples[1] = 16'b0000000000010100;
        samples[2] = 16'b0000000000100001;
        samples[3] = 16'b0000000010110001;
        samples[4] = 16'b1111111010101010;
        samples[5] = 16'b0000000100110100;
        samples[6] = 16'b0000000011111111;
        samples[7] = 16'b0000000011011100;
        samples[8] = 16'b1111101110100110;
        samples[9] = 16'b0000001111010100;
        samples[10] = 16'b0000000110100100;
        samples[11] = 16'b0000000101100000;
        samples[12] = 16'b1111111001001111;
        samples[13] = 16'b0000001100110101;
        samples[14] = 16'b1111111101111000;
        samples[15] = 16'b0000001001010011;
        samples[16] = 16'b0000000111110110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000100100111;
        samples[1] = 16'b0000000001111011;
        samples[2] = 16'b0000000010100100;
        samples[3] = 16'b0000000000101010;
        samples[4] = 16'b1111111101000000;
        samples[5] = 16'b0000000110110100;
        samples[6] = 16'b0000000100110100;
        samples[7] = 16'b0000000001010000;
        samples[8] = 16'b1111110011010010;
        samples[9] = 16'b0000001111101101;
        samples[10] = 16'b0000000101111111;
        samples[11] = 16'b0000000001101100;
        samples[12] = 16'b0000000101001101;
        samples[13] = 16'b0000001101001010;
        samples[14] = 16'b1111111001010101;
        samples[15] = 16'b0000001010110100;
        samples[16] = 16'b0000000111111001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110011000;
        samples[1] = 16'b0000000001111000;
        samples[2] = 16'b0000000010110100;
        samples[3] = 16'b0000000000101101;
        samples[4] = 16'b1111111111010011;
        samples[5] = 16'b0000000111100000;
        samples[6] = 16'b0000000100101110;
        samples[7] = 16'b0000000000100001;
        samples[8] = 16'b1111110011000010;
        samples[9] = 16'b0000001100100010;
        samples[10] = 16'b0000000110101011;
        samples[11] = 16'b0000000100011011;
        samples[12] = 16'b0000011000111001;
        samples[13] = 16'b1111110110000100;
        samples[14] = 16'b0000000001000000;
        samples[15] = 16'b0000001011100110;
        samples[16] = 16'b0000001000001100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000111000100;
        samples[1] = 16'b0000000001111111;
        samples[2] = 16'b0000000011100011;
        samples[3] = 16'b0000000001111000;
        samples[4] = 16'b0000000000101101;
        samples[5] = 16'b0000001000011110;
        samples[6] = 16'b0000000100110111;
        samples[7] = 16'b0000000000011110;
        samples[8] = 16'b1111110110110110;
        samples[9] = 16'b0000010001001110;
        samples[10] = 16'b0000000101010110;
        samples[11] = 16'b0000000100011011;
        samples[12] = 16'b0000000000111010;
        samples[13] = 16'b0000001001011101;
        samples[14] = 16'b1111111110010001;
        samples[15] = 16'b0000001100111000;
        samples[16] = 16'b0000001000101011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000110011011;
        samples[1] = 16'b0000000010101010;
        samples[2] = 16'b0000000011111000;
        samples[3] = 16'b0000000010001000;
        samples[4] = 16'b0000000010000010;
        samples[5] = 16'b0000001000001000;
        samples[6] = 16'b0000000011110101;
        samples[7] = 16'b0000000001001001;
        samples[8] = 16'b1111111001000011;
        samples[9] = 16'b0000010001011010;
        samples[10] = 16'b0000000010100100;
        samples[11] = 16'b0000000010101010;
        samples[12] = 16'b0000000111101100;
        samples[13] = 16'b0000010011100111;
        samples[14] = 16'b1111111110000101;
        samples[15] = 16'b0000001100110001;
        samples[16] = 16'b0000000111011010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101101001;
        samples[1] = 16'b0000000001110010;
        samples[2] = 16'b0000000011011100;
        samples[3] = 16'b0000000011000110;
        samples[4] = 16'b0000000001110101;
        samples[5] = 16'b0000000110110100;
        samples[6] = 16'b0000000010110100;
        samples[7] = 16'b0000000010011110;
        samples[8] = 16'b1111110110101101;
        samples[9] = 16'b0000010000101000;
        samples[10] = 16'b0000000011010110;
        samples[11] = 16'b0000000011011111;
        samples[12] = 16'b0000000101010110;
        samples[13] = 16'b0000000100100001;
        samples[14] = 16'b1111111110110111;
        samples[15] = 16'b0000001100100101;
        samples[16] = 16'b0000000110011110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101100011;
        samples[1] = 16'b0000000001000011;
        samples[2] = 16'b0000000100110001;
        samples[3] = 16'b0000000100000010;
        samples[4] = 16'b0000000010010100;
        samples[5] = 16'b0000000101110110;
        samples[6] = 16'b0000000011111111;
        samples[7] = 16'b0000000011010011;
        samples[8] = 16'b1111110101010101;
        samples[9] = 16'b0000010010101100;
        samples[10] = 16'b0000000101010000;
        samples[11] = 16'b0000000101001101;
        samples[12] = 16'b1111111101000000;
        samples[13] = 16'b0000001100000011;
        samples[14] = 16'b0000000000000010;
        samples[15] = 16'b0000001101011010;
        samples[16] = 16'b0000000111001101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101100011;
        samples[1] = 16'b0000000001011001;
        samples[2] = 16'b0000000101101100;
        samples[3] = 16'b0000000010010001;
        samples[4] = 16'b0000000011010110;
        samples[5] = 16'b0000000101000111;
        samples[6] = 16'b0000000100111010;
        samples[7] = 16'b0000000001011111;
        samples[8] = 16'b1111110111001111;
        samples[9] = 16'b0000010100000011;
        samples[10] = 16'b0000000100100111;
        samples[11] = 16'b0000000001100010;
        samples[12] = 16'b1111111101010110;
        samples[13] = 16'b0000011010001010;
        samples[14] = 16'b1111111111000000;
        samples[15] = 16'b0000001101101101;
        samples[16] = 16'b0000000111001010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101101100;
        samples[1] = 16'b0000000001001101;
        samples[2] = 16'b0000000101111001;
        samples[3] = 16'b0000000000010111;
        samples[4] = 16'b0000000011101001;
        samples[5] = 16'b0000000100110100;
        samples[6] = 16'b0000000011111000;
        samples[7] = 16'b0000000000110000;
        samples[8] = 16'b1111111000010100;
        samples[9] = 16'b0000001011111100;
        samples[10] = 16'b0000000110111101;
        samples[11] = 16'b0000000001110101;
        samples[12] = 16'b0000000110011011;
        samples[13] = 16'b0000000110100001;
        samples[14] = 16'b0000000001000000;
        samples[15] = 16'b0000001011111100;
        samples[16] = 16'b0000000110001000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000111000111;
        samples[1] = 16'b0000000001011111;
        samples[2] = 16'b0000000110101000;
        samples[3] = 16'b1111111110001110;
        samples[4] = 16'b0000000101011001;
        samples[5] = 16'b0000000101010000;
        samples[6] = 16'b0000000011100110;
        samples[7] = 16'b1111111111001100;
        samples[8] = 16'b1111110111000110;
        samples[9] = 16'b0000001100011000;
        samples[10] = 16'b0000001000011011;
        samples[11] = 16'b0000000010001110;
        samples[12] = 16'b0000000001101001;
        samples[13] = 16'b0000011000111100;
        samples[14] = 16'b0000000011101100;
        samples[15] = 16'b0000001011001010;
        samples[16] = 16'b0000000110000010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000101011001;
        samples[1] = 16'b0000000000111101;
        samples[2] = 16'b0000000101101100;
        samples[3] = 16'b1111111111011111;
        samples[4] = 16'b0000000100100111;
        samples[5] = 16'b0000000100001000;
        samples[6] = 16'b0000000010100001;
        samples[7] = 16'b0000000000001000;
        samples[8] = 16'b1111110111010101;
        samples[9] = 16'b0000001101001110;
        samples[10] = 16'b0000000110001000;
        samples[11] = 16'b0000000000110000;
        samples[12] = 16'b0000001000110111;
        samples[13] = 16'b0000000111001101;
        samples[14] = 16'b0000000101111100;
        samples[15] = 16'b0000001001101100;
        samples[16] = 16'b0000000100100001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000100000010;
        samples[1] = 16'b0000000000100001;
        samples[2] = 16'b0000000101100110;
        samples[3] = 16'b1111111111100101;
        samples[4] = 16'b0000000100100111;
        samples[5] = 16'b0000000011010110;
        samples[6] = 16'b0000000001101100;
        samples[7] = 16'b0000000000000010;
        samples[8] = 16'b1111111100011010;
        samples[9] = 16'b0000001101011010;
        samples[10] = 16'b0000000010101101;
        samples[11] = 16'b1111111110001000;
        samples[12] = 16'b0000000111011010;
        samples[13] = 16'b1111110011001011;
        samples[14] = 16'b0000000010001011;
        samples[15] = 16'b0000000111111111;
        samples[16] = 16'b0000000010101101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011100110;
        samples[1] = 16'b0000000000100001;
        samples[2] = 16'b0000000101100000;
        samples[3] = 16'b1111111111001100;
        samples[4] = 16'b0000000100100100;
        samples[5] = 16'b0000000010010001;
        samples[6] = 16'b0000000001010011;
        samples[7] = 16'b0000000000100100;
        samples[8] = 16'b1111110110110011;
        samples[9] = 16'b0000001110101110;
        samples[10] = 16'b0000000100100111;
        samples[11] = 16'b1111111111001001;
        samples[12] = 16'b0000001000111110;
        samples[13] = 16'b1111110001010010;
        samples[14] = 16'b0000000010010100;
        samples[15] = 16'b0000000110110001;
        samples[16] = 16'b0000000001110101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011100011;
        samples[1] = 16'b0000000000101101;
        samples[2] = 16'b0000000101010110;
        samples[3] = 16'b1111111111000000;
        samples[4] = 16'b0000000101110110;
        samples[5] = 16'b0000000001001001;
        samples[6] = 16'b0000000001010011;
        samples[7] = 16'b0000000000010001;
        samples[8] = 16'b1111111100110000;
        samples[9] = 16'b0000001110000011;
        samples[10] = 16'b0000000000100111;
        samples[11] = 16'b1111111100001000;
        samples[12] = 16'b0000010011100001;
        samples[13] = 16'b1111100110011111;
        samples[14] = 16'b1111111110010001;
        samples[15] = 16'b0000000101001010;
        samples[16] = 16'b0000000000100111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000010111101;
        samples[1] = 16'b0000000001000011;
        samples[2] = 16'b0000000100011011;
        samples[3] = 16'b1111111111000011;
        samples[4] = 16'b0000000101111001;
        samples[5] = 16'b1111111111011100;
        samples[6] = 16'b0000000000111010;
        samples[7] = 16'b0000000001001101;
        samples[8] = 16'b1111111011010101;
        samples[9] = 16'b0000001011010000;
        samples[10] = 16'b0000000010010100;
        samples[11] = 16'b1111111100100100;
        samples[12] = 16'b0000001111100000;
        samples[13] = 16'b1111110100111100;
        samples[14] = 16'b1111111110010001;
        samples[15] = 16'b0000000011011100;
        samples[16] = 16'b0000000000000010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011010011;
        samples[1] = 16'b0000000000100001;
        samples[2] = 16'b0000000011100110;
        samples[3] = 16'b1111111111101001;
        samples[4] = 16'b0000000110011110;
        samples[5] = 16'b1111111110000001;
        samples[6] = 16'b0000000000000101;
        samples[7] = 16'b0000000010011000;
        samples[8] = 16'b1111111001010010;
        samples[9] = 16'b0000001010110100;
        samples[10] = 16'b0000000010101010;
        samples[11] = 16'b1111111110111010;
        samples[12] = 16'b0000001101100011;
        samples[13] = 16'b0000001000001000;
        samples[14] = 16'b0000000000111010;
        samples[15] = 16'b0000000010011011;
        samples[16] = 16'b1111111110111101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000011000000;
        samples[1] = 16'b1111111111010110;
        samples[2] = 16'b0000000010111010;
        samples[3] = 16'b0000000001000000;
        samples[4] = 16'b0000000111101001;
        samples[5] = 16'b1111111100010111;
        samples[6] = 16'b1111111111010000;
        samples[7] = 16'b0000000011000011;
        samples[8] = 16'b0000000010010100;
        samples[9] = 16'b0000000110110100;
        samples[10] = 16'b1111111101100101;
        samples[11] = 16'b1111111111001100;
        samples[12] = 16'b0000000100111101;
        samples[13] = 16'b0000000011101111;
        samples[14] = 16'b0000000010001110;
        samples[15] = 16'b0000000000110111;
        samples[16] = 16'b1111111101000011;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000001100010;
        samples[1] = 16'b1111111111100010;
        samples[2] = 16'b0000000001110101;
        samples[3] = 16'b0000000001010110;
        samples[4] = 16'b0000000110101000;
        samples[5] = 16'b1111111011010101;
        samples[6] = 16'b1111111110101010;
        samples[7] = 16'b0000000011101111;
        samples[8] = 16'b1111111110001011;
        samples[9] = 16'b0000000100001000;
        samples[10] = 16'b0000000001101100;
        samples[11] = 16'b1111111110011110;
        samples[12] = 16'b1111111110001000;
        samples[13] = 16'b0000001011110110;
        samples[14] = 16'b0000000010011110;
        samples[15] = 16'b0000000000001000;
        samples[16] = 16'b1111111100010100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111111110101;
        samples[1] = 16'b1111111110110000;
        samples[2] = 16'b0000000000111010;
        samples[3] = 16'b0000000010100111;
        samples[4] = 16'b0000000110000101;
        samples[5] = 16'b1111111010100111;
        samples[6] = 16'b1111111101000011;
        samples[7] = 16'b0000000100011110;
        samples[8] = 16'b0000000101000100;
        samples[9] = 16'b0000000010100111;
        samples[10] = 16'b1111111010111001;
        samples[11] = 16'b1111111100001000;
        samples[12] = 16'b1111110010001101;
        samples[13] = 16'b0000001000011000;
        samples[14] = 16'b0000000001000011;
        samples[15] = 16'b1111111110011110;
        samples[16] = 16'b1111111010001110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000000100100;
        samples[1] = 16'b1111111110110000;
        samples[2] = 16'b0000000001011111;
        samples[3] = 16'b0000000000001110;
        samples[4] = 16'b0000000111011010;
        samples[5] = 16'b1111111011010101;
        samples[6] = 16'b1111111101011001;
        samples[7] = 16'b0000000001000011;
        samples[8] = 16'b0000001001110000;
        samples[9] = 16'b1111111110100100;
        samples[10] = 16'b1111111010010111;
        samples[11] = 16'b1111111011100101;
        samples[12] = 16'b1111110010111100;
        samples[13] = 16'b0000000001111000;
        samples[14] = 16'b0000000000100100;
        samples[15] = 16'b1111111101011001;
        samples[16] = 16'b1111111010010111;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b0000000000010001;
        samples[1] = 16'b1111111101100010;
        samples[2] = 16'b0000000000100111;
        samples[3] = 16'b0000000000000101;
        samples[4] = 16'b0000000110010010;
        samples[5] = 16'b1111111010100011;
        samples[6] = 16'b1111111101100101;
        samples[7] = 16'b0000000000001011;
        samples[8] = 16'b0000000110011110;
        samples[9] = 16'b1111111011101011;
        samples[10] = 16'b1111111101010110;
        samples[11] = 16'b1111111101011100;
        samples[12] = 16'b1111111011011001;
        samples[13] = 16'b0000000000110111;
        samples[14] = 16'b0000000010011110;
        samples[15] = 16'b1111111100100100;
        samples[16] = 16'b1111111010101010;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110010111;
        samples[1] = 16'b1111111100111101;
        samples[2] = 16'b0000000000110100;
        samples[3] = 16'b0000000001111111;
        samples[4] = 16'b0000000100101011;
        samples[5] = 16'b1111111010000100;
        samples[6] = 16'b1111111100110000;
        samples[7] = 16'b0000000010101101;
        samples[8] = 16'b0000000110110001;
        samples[9] = 16'b1111111100100111;
        samples[10] = 16'b1111111011000000;
        samples[11] = 16'b1111111101000000;
        samples[12] = 16'b1111110010010110;
        samples[13] = 16'b1111111101110101;
        samples[14] = 16'b1111111111100010;
        samples[15] = 16'b1111111011101110;
        samples[16] = 16'b1111111001101110;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110001110;
        samples[1] = 16'b1111111100011101;
        samples[2] = 16'b0000000001000011;
        samples[3] = 16'b0000000000101010;
        samples[4] = 16'b0000000100011011;
        samples[5] = 16'b1111111001011111;
        samples[6] = 16'b1111111101000110;
        samples[7] = 16'b0000000001011111;
        samples[8] = 16'b0000001000110111;
        samples[9] = 16'b1111111100101101;
        samples[10] = 16'b1111111000101101;
        samples[11] = 16'b1111111011011100;
        samples[12] = 16'b1111111001111000;
        samples[13] = 16'b1111110101110001;
        samples[14] = 16'b1111111110110000;
        samples[15] = 16'b1111111011100010;
        samples[16] = 16'b1111111001001100;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110000001;
        samples[1] = 16'b1111111100001011;
        samples[2] = 16'b0000000000011110;
        samples[3] = 16'b0000000000001110;
        samples[4] = 16'b0000000011011111;
        samples[5] = 16'b1111111000110110;
        samples[6] = 16'b1111111110100100;
        samples[7] = 16'b0000000000000010;
        samples[8] = 16'b0000000010000101;
        samples[9] = 16'b1111111101100101;
        samples[10] = 16'b1111111101010011;
        samples[11] = 16'b1111111100101010;
        samples[12] = 16'b1111111111011100;
        samples[13] = 16'b1111111001110001;
        samples[14] = 16'b0000000000011110;
        samples[15] = 16'b1111111011101110;
        samples[16] = 16'b1111111010010001;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111101001111;
        samples[1] = 16'b1111111010111001;
        samples[2] = 16'b1111111110110011;
        samples[3] = 16'b0000000001111011;
        samples[4] = 16'b0000000010001000;
        samples[5] = 16'b1111111000010001;
        samples[6] = 16'b1111111101101100;
        samples[7] = 16'b0000000000101101;
        samples[8] = 16'b0000000000110000;
        samples[9] = 16'b1111111110011010;
        samples[10] = 16'b1111111101011111;
        samples[11] = 16'b1111111100101101;
        samples[12] = 16'b1111110110111111;
        samples[13] = 16'b1111110000000000;
        samples[14] = 16'b0000000001111011;
        samples[15] = 16'b1111111011011001;
        samples[16] = 16'b1111111001111000;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110010100;
        samples[1] = 16'b1111111011101110;
        samples[2] = 16'b1111111110001110;
        samples[3] = 16'b1111111110111101;
        samples[4] = 16'b0000000011111000;
        samples[5] = 16'b1111111001001001;
        samples[6] = 16'b1111111100011010;
        samples[7] = 16'b1111111101101000;
        samples[8] = 16'b0000000011000110;
        samples[9] = 16'b1111111101000110;
        samples[10] = 16'b1111111010101101;
        samples[11] = 16'b1111111011010010;
        samples[12] = 16'b1111111001011100;
        samples[13] = 16'b1111110101111110;
        samples[14] = 16'b0000000100100100;
        samples[15] = 16'b1111111010000100;
        samples[16] = 16'b1111111001100101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)

        en = 1;
        samples[0] = 16'b1111111110101010;
        samples[1] = 16'b1111111011010101;
        samples[2] = 16'b1111111100110000;
        samples[3] = 16'b1111111110100001;
        samples[4] = 16'b0000000011101001;
        samples[5] = 16'b1111111000111001;
        samples[6] = 16'b1111111011100101;
        samples[7] = 16'b1111111100111101;
        samples[8] = 16'b0000000010011110;
        samples[9] = 16'b1111111100111010;
        samples[10] = 16'b1111111011000011;
        samples[11] = 16'b1111111100010001;
        samples[12] = 16'b1111111111000110;
        samples[13] = 16'b1111101101111101;
        samples[14] = 16'b0000000100111010;
        samples[15] = 16'b1111111001101011;
        samples[16] = 16'b1111111001010101;
       # (0.5 + 0.5)
        en = 0;
        # (3906.25 - 0.5- 0.5)
        $vcdplusfile("tb_ma_encoder_mapped.vpd");
        $vcdpluson;

        $dumpfile("ma_encoder_mapped.dump");
        $dumpvars(0,tb_ma_encoder_mapped);
        $dumpon;
        en = 1;
        samples[0] = 16'b1111111101001111;
        samples[1] = 16'b1111111010100111;
        samples[2] = 16'b1111111100101101;
        samples[3] = 16'b0000000000000010;
        samples[4] = 16'b0000000010011011;
        samples[5] = 16'b1111111000010100;
        samples[6] = 16'b1111111011010010;
        samples[7] = 16'b1111111110010001;
        samples[8] = 16'b0000000011111000;
        samples[9] = 16'b1111111100011101;
        samples[10] = 16'b1111111001111000;
        samples[11] = 16'b1111111011111110;
        samples[12] = 16'b1111111000010001;
        samples[13] = 16'b1111110001000010;
        samples[14] = 16'b0000000100100001;
        samples[15] = 16'b1111111001001001;
        samples[16] = 16'b1111111000110011;
       # (0.5 + 0.5)
        en = 0;

        wait (u_ma_encoder.done == 1);
        $dumpoff;
        # 2
        $finish;
    end
endmodule